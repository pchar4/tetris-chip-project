magic
tech scmos
timestamp 1711653199
<< metal1 >>
rect 14 3307 3458 3327
rect 38 3283 3434 3303
rect 14 3267 3458 3273
rect 196 3213 221 3216
rect 258 3213 284 3216
rect 410 3213 444 3216
rect 492 3213 517 3216
rect 604 3213 629 3216
rect 660 3213 701 3216
rect 722 3213 765 3216
rect 802 3213 828 3216
rect 900 3213 925 3216
rect 970 3213 996 3216
rect 1044 3213 1069 3216
rect 1180 3213 1189 3216
rect 1258 3213 1276 3216
rect 1316 3213 1333 3216
rect 1420 3213 1445 3216
rect 1476 3213 1485 3216
rect 1556 3213 1581 3216
rect 1612 3213 1621 3216
rect 1628 3213 1637 3216
rect 1684 3213 1709 3216
rect 1788 3213 1813 3216
rect 1844 3213 1853 3216
rect 1860 3213 1877 3216
rect 1916 3213 1941 3216
rect 1972 3213 1981 3216
rect 2020 3213 2045 3216
rect 2116 3213 2141 3216
rect 2172 3213 2181 3216
rect 2364 3213 2389 3216
rect 2420 3213 2429 3216
rect 2908 3213 2917 3216
rect 2996 3213 3021 3216
rect 3052 3213 3077 3216
rect 3172 3213 3181 3216
rect 3228 3213 3253 3216
rect 3284 3213 3293 3216
rect 674 3203 700 3206
rect 746 3203 772 3206
rect 1482 3205 1485 3213
rect 1618 3205 1621 3213
rect 1850 3205 1853 3213
rect 2178 3205 2181 3213
rect 2426 3205 2429 3213
rect 2914 3206 2917 3213
rect 2914 3203 2924 3206
rect 38 3167 3434 3173
rect 1106 3143 1116 3146
rect 1266 3143 1284 3146
rect 1386 3143 1396 3146
rect 1850 3143 1860 3146
rect 2122 3143 2132 3146
rect 2146 3143 2157 3146
rect 2298 3143 2308 3146
rect 3138 3143 3148 3146
rect 3170 3143 3188 3146
rect 3314 3143 3332 3146
rect 2154 3136 2157 3143
rect 234 3133 252 3136
rect 276 3133 301 3136
rect 442 3133 452 3136
rect 914 3133 924 3136
rect 1018 3133 1044 3136
rect 1106 3133 1124 3136
rect 1138 3133 1164 3136
rect 1234 3133 1252 3136
rect 1282 3133 1292 3136
rect 1378 3133 1404 3136
rect 1410 3133 1428 3136
rect 1434 3133 1468 3136
rect 1498 3133 1508 3136
rect 1522 3133 1540 3136
rect 1564 3133 1573 3136
rect 1628 3133 1661 3136
rect 1740 3133 1757 3136
rect 1762 3133 1788 3136
rect 234 3126 237 3133
rect 1498 3126 1501 3133
rect 1810 3126 1813 3135
rect 1868 3133 1909 3136
rect 1940 3133 1949 3136
rect 1988 3133 2013 3136
rect 2140 3133 2149 3136
rect 2154 3133 2164 3136
rect 2202 3133 2212 3136
rect 2292 3133 2301 3136
rect 2420 3133 2437 3136
rect 2762 3133 2780 3136
rect 2986 3133 3012 3136
rect 3026 3133 3052 3136
rect 3058 3133 3068 3136
rect 3106 3133 3116 3136
rect 3130 3133 3156 3136
rect 3178 3133 3196 3136
rect 3314 3133 3340 3136
rect 196 3123 212 3126
rect 226 3123 237 3126
rect 340 3123 365 3126
rect 402 3123 436 3126
rect 450 3123 460 3126
rect 474 3123 500 3126
rect 514 3123 532 3126
rect 604 3123 629 3126
rect 660 3123 669 3126
rect 716 3123 741 3126
rect 772 3123 781 3126
rect 796 3123 805 3126
rect 844 3123 869 3126
rect 906 3123 932 3126
rect 978 3123 988 3126
rect 1010 3123 1052 3126
rect 1066 3123 1084 3126
rect 1132 3123 1172 3126
rect 1260 3123 1277 3126
rect 1300 3123 1316 3126
rect 1330 3123 1356 3126
rect 1436 3123 1469 3126
rect 1490 3123 1501 3126
rect 1692 3123 1708 3126
rect 1810 3123 1821 3126
rect 1924 3123 1933 3126
rect 1948 3123 1964 3126
rect 2002 3123 2044 3126
rect 2148 3123 2172 3126
rect 2268 3123 2277 3126
rect 2300 3123 2309 3126
rect 2330 3123 2372 3126
rect 2476 3123 2485 3126
rect 2562 3123 2580 3126
rect 2642 3123 2652 3126
rect 2690 3123 2708 3126
rect 2820 3123 2829 3126
rect 2924 3123 2949 3126
rect 3020 3123 3037 3126
rect 3066 3123 3076 3126
rect 3082 3123 3124 3126
rect 3164 3123 3181 3126
rect 3228 3123 3276 3126
rect 3290 3123 3308 3126
rect 228 3113 237 3116
rect 276 3113 301 3116
rect 468 3113 477 3116
rect 514 3115 517 3123
rect 540 3113 565 3116
rect 1004 3113 1021 3116
rect 1332 3113 1341 3116
rect 2060 3113 2085 3116
rect 2188 3113 2197 3116
rect 3132 3113 3141 3116
rect 2082 3106 2085 3113
rect 2082 3103 2101 3106
rect 90 3083 173 3086
rect 14 3067 3458 3073
rect 2154 3033 2188 3036
rect 2418 3033 2460 3036
rect 356 3023 381 3026
rect 588 3023 613 3026
rect 660 3023 677 3026
rect 3108 3023 3117 3026
rect 3242 3016 3245 3025
rect 116 3013 133 3016
rect 172 3013 197 3016
rect 308 3013 340 3016
rect 404 3013 413 3016
rect 514 3013 540 3016
rect 602 3013 620 3016
rect 812 3013 828 3016
rect 876 3013 892 3016
rect 898 3013 932 3016
rect 954 3013 972 3016
rect 194 3005 197 3013
rect 1034 3006 1037 3014
rect 1090 3013 1108 3016
rect 1164 3013 1204 3016
rect 1234 3013 1244 3016
rect 1268 3013 1293 3016
rect 1362 3013 1380 3016
rect 1394 3013 1405 3016
rect 1426 3013 1469 3016
rect 1516 3013 1525 3016
rect 1532 3013 1541 3016
rect 1762 3013 1772 3016
rect 1802 3013 1836 3016
rect 1866 3013 1876 3016
rect 1948 3013 1965 3016
rect 2060 3013 2069 3016
rect 2076 3013 2092 3016
rect 2130 3013 2140 3016
rect 2228 3013 2237 3016
rect 2244 3013 2269 3016
rect 252 3003 285 3006
rect 300 3003 309 3006
rect 356 3003 365 3006
rect 396 3003 405 3006
rect 594 3003 612 3006
rect 626 3003 636 3006
rect 762 3003 788 3006
rect 810 3003 820 3006
rect 834 3003 852 3006
rect 874 3003 884 3006
rect 1034 3003 1052 3006
rect 1090 3003 1100 3006
rect 1146 3003 1156 3006
rect 1162 3003 1196 3006
rect 1250 3003 1260 3006
rect 1266 3003 1292 3006
rect 1402 3005 1405 3013
rect 1428 3003 1437 3006
rect 1612 3003 1628 3006
rect 1684 3003 1700 3006
rect 1724 3003 1733 3006
rect 1754 3003 1764 3006
rect 1802 3003 1828 3006
rect 2010 3003 2036 3006
rect 2082 3003 2100 3006
rect 2202 3003 2220 3006
rect 2266 3005 2269 3013
rect 2306 3006 2309 3014
rect 2364 3013 2373 3016
rect 2394 3013 2412 3016
rect 2500 3013 2524 3016
rect 2562 3013 2613 3016
rect 2682 3013 2716 3016
rect 2844 3013 2869 3016
rect 2900 3013 2909 3016
rect 2946 3013 2964 3016
rect 2978 3013 2988 3016
rect 3042 3013 3085 3016
rect 3138 3013 3148 3016
rect 3154 3013 3196 3016
rect 3242 3013 3253 3016
rect 3340 3013 3357 3016
rect 2906 3006 2909 3013
rect 2282 3003 2292 3006
rect 2306 3003 2341 3006
rect 2362 3003 2380 3006
rect 2474 3003 2484 3006
rect 2548 3003 2557 3006
rect 2578 3003 2612 3006
rect 2626 3003 2636 3006
rect 2650 3003 2660 3006
rect 2796 3003 2805 3006
rect 2906 3003 2916 3006
rect 2970 3003 2980 3006
rect 3058 3003 3068 3006
rect 3082 3003 3092 3006
rect 3170 3003 3188 3006
rect 3250 3005 3253 3013
rect 226 2993 244 2996
rect 258 2993 292 2996
rect 362 2993 388 2996
rect 834 2993 837 3003
rect 1458 2993 1484 2996
rect 1586 2993 1604 2996
rect 1666 2993 1676 2996
rect 1730 2993 1740 2996
rect 2082 2983 2085 3003
rect 2970 2983 2973 3003
rect 38 2967 3434 2973
rect 1226 2936 1229 2946
rect 1282 2943 1292 2946
rect 514 2933 524 2936
rect 538 2933 556 2936
rect 634 2933 644 2936
rect 658 2933 684 2936
rect 716 2933 725 2936
rect 930 2933 940 2936
rect 1026 2933 1044 2936
rect 1132 2933 1165 2936
rect 1226 2933 1236 2936
rect 2018 2933 2036 2936
rect 2076 2933 2093 2936
rect 2332 2933 2349 2936
rect 2634 2933 2644 2936
rect 2690 2933 2708 2936
rect 3138 2933 3148 2936
rect 3154 2933 3164 2936
rect 3234 2933 3252 2936
rect 3276 2933 3301 2936
rect 514 2926 517 2933
rect 634 2926 637 2933
rect 116 2923 141 2926
rect 212 2923 228 2926
rect 356 2923 365 2926
rect 506 2923 517 2926
rect 554 2923 564 2926
rect 626 2923 637 2926
rect 692 2923 701 2926
rect 762 2923 772 2926
rect 778 2923 812 2926
rect 866 2923 876 2926
rect 890 2923 941 2926
rect 1034 2923 1076 2926
rect 1106 2923 1116 2926
rect 1218 2923 1244 2926
rect 1276 2923 1285 2926
rect 1426 2923 1444 2926
rect 1596 2923 1621 2926
rect 1658 2923 1668 2926
rect 1732 2923 1741 2926
rect 1836 2923 1861 2926
rect 1908 2923 1925 2926
rect 244 2913 261 2916
rect 580 2913 597 2916
rect 732 2913 741 2916
rect 828 2913 837 2916
rect 956 2913 973 2916
rect 988 2913 997 2916
rect 1212 2913 1229 2916
rect 1340 2913 1365 2916
rect 1420 2913 1429 2916
rect 1460 2913 1469 2916
rect 1508 2913 1517 2916
rect 1684 2913 1693 2916
rect 1948 2913 1957 2916
rect 2090 2906 2093 2933
rect 2130 2923 2157 2926
rect 2196 2923 2213 2926
rect 2346 2925 2349 2933
rect 2500 2923 2509 2926
rect 2610 2923 2628 2926
rect 2634 2923 2652 2926
rect 2716 2923 2725 2926
rect 2924 2923 2941 2926
rect 3076 2923 3101 2926
rect 3236 2923 3245 2926
rect 2210 2906 2213 2923
rect 2276 2913 2285 2916
rect 2300 2913 2317 2916
rect 2418 2913 2436 2916
rect 2986 2913 3004 2916
rect 3036 2913 3045 2916
rect 3090 2913 3108 2916
rect 730 2903 748 2906
rect 962 2903 980 2906
rect 1186 2903 1204 2906
rect 1314 2903 1332 2906
rect 1466 2903 1500 2906
rect 1946 2903 1964 2906
rect 2090 2903 2116 2906
rect 2210 2903 2236 2906
rect 2274 2903 2292 2906
rect 2394 2903 2404 2906
rect 2994 2903 3020 2906
rect 3034 2903 3052 2906
rect 3106 2903 3124 2906
rect 14 2867 3458 2873
rect 3068 2823 3085 2826
rect 3082 2816 3085 2823
rect 148 2813 173 2816
rect 284 2813 325 2816
rect 386 2813 404 2816
rect 436 2813 453 2816
rect 458 2813 468 2816
rect 594 2813 604 2816
rect 636 2813 661 2816
rect 714 2813 732 2816
rect 778 2813 796 2816
rect 828 2813 853 2816
rect 892 2813 909 2816
rect 922 2806 925 2814
rect 956 2813 989 2816
rect 1028 2813 1045 2816
rect 1090 2813 1125 2816
rect 1130 2813 1172 2816
rect 1244 2813 1261 2816
rect 1436 2813 1453 2816
rect 1612 2813 1621 2816
rect 1810 2813 1836 2816
rect 1932 2813 1957 2816
rect 1996 2813 2021 2816
rect 2100 2813 2125 2816
rect 2196 2813 2213 2816
rect 2396 2813 2421 2816
rect 2676 2813 2701 2816
rect 3002 2813 3020 2816
rect 3026 2813 3060 2816
rect 3082 2813 3093 2816
rect 3114 2813 3132 2816
rect 3284 2813 3293 2816
rect 3308 2813 3317 2816
rect 3332 2813 3356 2816
rect 3388 2813 3397 2816
rect 140 2803 189 2806
rect 290 2803 340 2806
rect 356 2803 373 2806
rect 402 2803 412 2806
rect 434 2803 476 2806
rect 570 2803 612 2806
rect 634 2803 660 2806
rect 714 2803 724 2806
rect 762 2803 804 2806
rect 826 2803 868 2806
rect 890 2803 925 2806
rect 1122 2803 1164 2806
rect 1196 2803 1236 2806
rect 1386 2803 1412 2806
rect 1858 2803 1868 2806
rect 1890 2803 1908 2806
rect 2458 2803 2468 2806
rect 2602 2803 2612 2806
rect 2668 2803 2677 2806
rect 3004 2803 3012 2806
rect 3090 2805 3093 2813
rect 3116 2803 3124 2806
rect 3188 2803 3197 2806
rect 3212 2803 3221 2806
rect 2458 2783 2461 2803
rect 3306 2793 3316 2796
rect 38 2767 3434 2773
rect 202 2726 205 2735
rect 442 2726 445 2735
rect 116 2723 141 2726
rect 172 2723 205 2726
rect 212 2723 228 2726
rect 332 2723 357 2726
rect 388 2723 397 2726
rect 402 2723 420 2726
rect 434 2723 445 2726
rect 466 2726 469 2735
rect 474 2733 508 2736
rect 562 2733 572 2736
rect 698 2733 740 2736
rect 780 2733 797 2736
rect 858 2733 885 2736
rect 914 2733 924 2736
rect 954 2733 964 2736
rect 1098 2733 1124 2736
rect 1204 2733 1229 2736
rect 562 2726 565 2733
rect 466 2723 477 2726
rect 554 2723 565 2726
rect 610 2723 628 2726
rect 658 2723 668 2726
rect 748 2723 757 2726
rect 468 2713 493 2716
rect 794 2706 797 2733
rect 1250 2726 1253 2735
rect 1266 2733 1300 2736
rect 1322 2733 1348 2736
rect 1946 2733 1972 2736
rect 2148 2733 2156 2736
rect 2282 2733 2324 2736
rect 2346 2733 2372 2736
rect 2530 2733 2556 2736
rect 2908 2733 2933 2736
rect 3018 2733 3028 2736
rect 3250 2733 3260 2736
rect 842 2723 852 2726
rect 866 2723 908 2726
rect 946 2723 956 2726
rect 1058 2723 1076 2726
rect 1090 2723 1141 2726
rect 1212 2723 1253 2726
rect 1260 2723 1285 2726
rect 1372 2723 1381 2726
rect 1652 2723 1661 2726
rect 1858 2723 1884 2726
rect 1906 2723 1924 2726
rect 1996 2723 2021 2726
rect 2060 2723 2077 2726
rect 2122 2723 2132 2726
rect 2164 2723 2181 2726
rect 2220 2723 2245 2726
rect 2306 2723 2316 2726
rect 2348 2723 2357 2726
rect 2396 2723 2421 2726
rect 2580 2723 2589 2726
rect 2636 2723 2661 2726
rect 2890 2723 2901 2726
rect 2916 2723 2948 2726
rect 3092 2723 3117 2726
rect 3282 2723 3300 2726
rect 3348 2724 3364 2727
rect 2890 2716 2893 2723
rect 802 2713 812 2716
rect 836 2713 845 2716
rect 860 2713 893 2716
rect 2876 2713 2893 2716
rect 3004 2713 3013 2716
rect 3380 2713 3389 2716
rect 794 2703 828 2706
rect 1154 2703 1180 2706
rect 3362 2703 3372 2706
rect 14 2667 3458 2673
rect 1082 2633 1116 2636
rect 1178 2633 1204 2636
rect 388 2623 405 2626
rect 556 2623 565 2626
rect 588 2623 605 2626
rect 620 2623 629 2626
rect 700 2623 717 2626
rect 116 2613 133 2616
rect 172 2613 197 2616
rect 244 2613 261 2616
rect 300 2613 325 2616
rect 444 2613 469 2616
rect 500 2613 517 2616
rect 524 2613 540 2616
rect 570 2613 580 2616
rect 586 2613 612 2616
rect 634 2613 652 2616
rect 674 2613 684 2616
rect 698 2613 732 2616
rect 764 2613 781 2616
rect 178 2603 212 2606
rect 218 2603 236 2606
rect 388 2603 397 2606
rect 514 2605 517 2613
rect 786 2606 789 2614
rect 874 2613 900 2616
rect 1082 2606 1085 2633
rect 1162 2623 1188 2626
rect 2962 2616 2965 2625
rect 1130 2613 1140 2616
rect 1146 2613 1156 2616
rect 1250 2613 1276 2616
rect 1306 2613 1316 2616
rect 1524 2613 1549 2616
rect 1580 2613 1613 2616
rect 1740 2613 1765 2616
rect 1796 2613 1813 2616
rect 1964 2613 1997 2616
rect 2188 2613 2221 2616
rect 2260 2613 2285 2616
rect 2364 2613 2389 2616
rect 2580 2613 2597 2616
rect 2676 2613 2709 2616
rect 2724 2613 2741 2616
rect 2922 2613 2948 2616
rect 2962 2613 2980 2616
rect 3018 2613 3028 2616
rect 562 2603 572 2606
rect 706 2603 724 2606
rect 778 2603 789 2606
rect 812 2603 829 2606
rect 858 2603 892 2606
rect 1068 2603 1085 2606
rect 1228 2603 1261 2606
rect 1300 2603 1308 2606
rect 1610 2605 1613 2613
rect 1636 2603 1652 2606
rect 1676 2603 1701 2606
rect 1810 2605 1813 2613
rect 1860 2603 1869 2606
rect 1994 2605 1997 2613
rect 3050 2606 3053 2614
rect 3068 2613 3084 2616
rect 3146 2606 3149 2614
rect 3180 2613 3205 2616
rect 3332 2613 3349 2616
rect 2010 2603 2020 2606
rect 2076 2603 2124 2606
rect 2146 2603 2164 2606
rect 2716 2603 2741 2606
rect 2746 2603 2756 2606
rect 2772 2603 2781 2606
rect 2842 2603 2868 2606
rect 2930 2603 2940 2606
rect 2994 2603 3036 2606
rect 3050 2603 3060 2606
rect 3074 2603 3092 2606
rect 3114 2603 3149 2606
rect 3178 2603 3188 2606
rect 3282 2603 3308 2606
rect 3330 2603 3372 2606
rect 562 2593 565 2603
rect 778 2593 781 2603
rect 1042 2593 1060 2596
rect 38 2567 3434 2573
rect 1130 2543 1156 2546
rect 1482 2543 1492 2546
rect 1602 2543 1636 2546
rect 1794 2543 1804 2546
rect 178 2533 205 2536
rect 228 2533 245 2536
rect 356 2533 373 2536
rect 506 2533 524 2536
rect 116 2523 133 2526
rect 172 2523 197 2526
rect 202 2525 205 2533
rect 674 2526 677 2535
rect 890 2526 893 2535
rect 1082 2533 1092 2536
rect 1124 2533 1141 2536
rect 1164 2533 1173 2536
rect 1370 2526 1373 2535
rect 1458 2533 1476 2536
rect 1500 2533 1525 2536
rect 1554 2526 1557 2535
rect 1594 2533 1644 2536
rect 1690 2533 1700 2536
rect 1706 2533 1748 2536
rect 1788 2533 1805 2536
rect 1812 2533 1845 2536
rect 2106 2533 2124 2536
rect 2428 2533 2437 2536
rect 2732 2533 2741 2536
rect 2764 2533 2781 2536
rect 3090 2533 3108 2536
rect 3178 2533 3196 2536
rect 3236 2533 3245 2536
rect 3300 2533 3309 2536
rect 1690 2526 1693 2533
rect 276 2523 285 2526
rect 340 2523 349 2526
rect 444 2523 469 2526
rect 500 2523 509 2526
rect 532 2523 541 2526
rect 588 2523 605 2526
rect 644 2523 677 2526
rect 684 2523 700 2526
rect 714 2523 732 2526
rect 812 2523 837 2526
rect 868 2523 893 2526
rect 900 2523 916 2526
rect 930 2523 948 2526
rect 970 2523 1004 2526
rect 1082 2523 1100 2526
rect 1194 2523 1204 2526
rect 1292 2523 1317 2526
rect 1348 2523 1373 2526
rect 1380 2523 1396 2526
rect 1418 2523 1436 2526
rect 1484 2523 1493 2526
rect 1514 2523 1540 2526
rect 1554 2523 1565 2526
rect 1658 2523 1668 2526
rect 1682 2523 1693 2526
rect 1708 2523 1749 2526
rect 1988 2523 2005 2526
rect 2044 2523 2069 2526
rect 2212 2523 2237 2526
rect 2324 2523 2349 2526
rect 2476 2523 2501 2526
rect 2532 2523 2541 2526
rect 2580 2523 2605 2526
rect 2636 2523 2645 2526
rect 2708 2523 2740 2526
rect 2836 2523 2861 2526
rect 2930 2523 2948 2526
rect 3028 2523 3053 2526
rect 714 2515 717 2523
rect 930 2515 933 2523
rect 1412 2513 1421 2516
rect 1452 2513 1461 2516
rect 2428 2513 2437 2516
rect 3090 2483 3093 2533
rect 3162 2523 3204 2526
rect 3164 2513 3173 2516
rect 3236 2513 3245 2516
rect 3322 2503 3325 2515
rect 3354 2503 3372 2506
rect 14 2467 3458 2473
rect 242 2453 285 2456
rect 3298 2433 3325 2436
rect 1666 2423 1676 2426
rect 2300 2423 2317 2426
rect 2388 2423 2397 2426
rect 2468 2423 2485 2426
rect 2612 2423 2621 2426
rect 3298 2423 3316 2426
rect 1666 2416 1669 2423
rect 364 2413 373 2416
rect 420 2413 437 2416
rect 484 2413 501 2416
rect 604 2413 621 2416
rect 812 2413 829 2416
rect 868 2413 893 2416
rect 1060 2413 1077 2416
rect 1156 2413 1165 2416
rect 1308 2413 1317 2416
rect 1346 2413 1396 2416
rect 1410 2413 1421 2416
rect 1588 2413 1597 2416
rect 1660 2413 1669 2416
rect 1706 2413 1716 2416
rect 1860 2413 1877 2416
rect 1956 2413 1981 2416
rect 2060 2413 2085 2416
rect 2164 2413 2181 2416
rect 2226 2413 2252 2416
rect 2266 2413 2277 2416
rect 2322 2413 2332 2416
rect 2362 2413 2372 2416
rect 2524 2413 2549 2416
rect 2586 2413 2596 2416
rect 2668 2413 2693 2416
rect 2724 2413 2741 2416
rect 2762 2413 2780 2416
rect 3050 2413 3076 2416
rect 3090 2413 3109 2416
rect 3130 2413 3156 2416
rect 3170 2413 3189 2416
rect 3244 2413 3253 2416
rect 3322 2415 3325 2433
rect 3372 2413 3381 2416
rect 700 2403 717 2406
rect 948 2403 965 2406
rect 1108 2403 1125 2406
rect 1154 2403 1196 2406
rect 1258 2403 1284 2406
rect 1306 2403 1316 2406
rect 1340 2403 1373 2406
rect 1378 2403 1388 2406
rect 1410 2405 1413 2413
rect 1468 2403 1477 2406
rect 1628 2403 1637 2406
rect 1722 2403 1732 2406
rect 1866 2403 1892 2406
rect 2266 2405 2269 2413
rect 2306 2403 2324 2406
rect 2348 2403 2357 2406
rect 2402 2403 2412 2406
rect 2730 2403 2740 2406
rect 2986 2403 2996 2406
rect 3090 2405 3093 2413
rect 3098 2403 3108 2406
rect 3170 2405 3173 2413
rect 3178 2403 3196 2406
rect 3258 2403 3276 2406
rect 1378 2396 1381 2403
rect 666 2393 692 2396
rect 930 2393 940 2396
rect 1362 2393 1381 2396
rect 114 2383 173 2386
rect 2730 2383 2733 2403
rect 3250 2393 3268 2396
rect 38 2367 3434 2373
rect 618 2333 628 2336
rect 898 2333 924 2336
rect 1258 2333 1276 2336
rect 1300 2333 1317 2336
rect 1618 2333 1628 2336
rect 1690 2333 1716 2336
rect 1874 2333 1908 2336
rect 1986 2333 2004 2336
rect 2034 2333 2068 2336
rect 2322 2333 2372 2336
rect 2428 2333 2437 2336
rect 2770 2333 2796 2336
rect 2828 2333 2837 2336
rect 2874 2333 2916 2336
rect 116 2323 125 2326
rect 172 2323 181 2326
rect 220 2323 245 2326
rect 276 2323 285 2326
rect 332 2323 357 2326
rect 436 2323 453 2326
rect 492 2323 509 2326
rect 618 2303 621 2333
rect 1690 2326 1693 2333
rect 836 2323 861 2326
rect 922 2323 932 2326
rect 1068 2323 1093 2326
rect 1180 2323 1205 2326
rect 1380 2323 1405 2326
rect 1442 2323 1460 2326
rect 1540 2323 1565 2326
rect 1610 2323 1636 2326
rect 1650 2323 1668 2326
rect 1682 2323 1693 2326
rect 1812 2323 1837 2326
rect 1874 2323 1916 2326
rect 1986 2323 2012 2326
rect 2026 2323 2076 2326
rect 2098 2323 2116 2326
rect 2210 2323 2269 2326
rect 1300 2313 1325 2316
rect 1476 2313 1485 2316
rect 2028 2313 2053 2316
rect 2258 2313 2276 2316
rect 2282 2306 2285 2325
rect 2306 2323 2316 2326
rect 2322 2323 2325 2333
rect 3114 2326 3117 2334
rect 3164 2333 3189 2336
rect 3290 2333 3316 2336
rect 3330 2333 3340 2336
rect 3354 2333 3364 2336
rect 2354 2323 2380 2326
rect 2492 2323 2517 2326
rect 2620 2323 2645 2326
rect 2676 2323 2693 2326
rect 2730 2323 2773 2326
rect 2778 2323 2804 2326
rect 3028 2323 3053 2326
rect 3084 2323 3117 2326
rect 3124 2323 3133 2326
rect 3138 2323 3148 2326
rect 3298 2323 3324 2326
rect 3338 2323 3348 2326
rect 3362 2323 3372 2326
rect 2770 2316 2773 2323
rect 2770 2313 2789 2316
rect 3164 2313 3189 2316
rect 3212 2313 3221 2316
rect 3332 2313 3341 2316
rect 2258 2303 2285 2306
rect 3178 2303 3228 2306
rect 3250 2303 3260 2306
rect 14 2267 3458 2273
rect 1202 2233 1244 2236
rect 1378 2233 1397 2236
rect 1994 2233 2021 2236
rect 2266 2233 2285 2236
rect 2306 2233 2317 2236
rect 2338 2233 2372 2236
rect 2394 2233 2404 2236
rect 2418 2233 2444 2236
rect 364 2223 381 2226
rect 508 2223 525 2226
rect 956 2223 997 2226
rect 1028 2223 1053 2226
rect 1138 2216 1141 2225
rect 1228 2223 1237 2226
rect 1252 2223 1277 2226
rect 1378 2216 1381 2233
rect 116 2213 133 2216
rect 234 2213 244 2216
rect 290 2213 332 2216
rect 338 2213 348 2216
rect 370 2213 412 2216
rect 586 2213 636 2216
rect 748 2213 765 2216
rect 868 2213 877 2216
rect 922 2213 940 2216
rect 970 2213 1012 2216
rect 1026 2213 1077 2216
rect 762 2206 765 2213
rect 186 2203 204 2206
rect 282 2203 324 2206
rect 394 2203 404 2206
rect 444 2203 453 2206
rect 458 2203 484 2206
rect 588 2203 605 2206
rect 642 2203 652 2206
rect 762 2203 780 2206
rect 802 2203 860 2206
rect 866 2203 876 2206
rect 962 2203 1004 2206
rect 1026 2205 1029 2213
rect 1034 2203 1084 2206
rect 1090 2196 1093 2214
rect 1106 2213 1124 2216
rect 1138 2213 1149 2216
rect 1156 2213 1181 2216
rect 1194 2206 1197 2214
rect 1298 2213 1308 2216
rect 1330 2213 1381 2216
rect 1394 2215 1397 2233
rect 1684 2223 1725 2226
rect 1756 2223 1765 2226
rect 1804 2223 1813 2226
rect 2002 2223 2012 2226
rect 1458 2206 1461 2214
rect 1516 2213 1525 2216
rect 1580 2213 1597 2216
rect 1642 2213 1668 2216
rect 1682 2213 1740 2216
rect 1754 2213 1765 2216
rect 1778 2213 1788 2216
rect 1802 2213 1820 2216
rect 1850 2213 1867 2216
rect 1898 2213 1925 2216
rect 1988 2213 2005 2216
rect 2018 2215 2021 2233
rect 2036 2223 2045 2226
rect 2228 2223 2237 2226
rect 2258 2223 2276 2226
rect 2282 2215 2285 2233
rect 2314 2215 2317 2233
rect 2338 2223 2356 2226
rect 2418 2223 2428 2226
rect 2458 2213 2492 2216
rect 1098 2203 1116 2206
rect 1162 2203 1188 2206
rect 1194 2203 1221 2206
rect 1258 2203 1300 2206
rect 1418 2203 1452 2206
rect 1458 2203 1508 2206
rect 1514 2203 1524 2206
rect 1538 2203 1572 2206
rect 1586 2203 1660 2206
rect 1682 2205 1685 2213
rect 1762 2206 1765 2213
rect 1850 2206 1853 2213
rect 1922 2206 1925 2213
rect 2514 2206 2517 2214
rect 2540 2213 2549 2216
rect 2588 2213 2613 2216
rect 2684 2213 2701 2216
rect 2738 2206 2741 2226
rect 3218 2216 3221 2225
rect 2802 2213 2820 2216
rect 2900 2213 2909 2216
rect 3004 2213 3029 2216
rect 3116 2213 3125 2216
rect 3178 2213 3204 2216
rect 3218 2213 3229 2216
rect 3244 2213 3308 2216
rect 3330 2213 3340 2216
rect 1762 2203 1780 2206
rect 1842 2203 1853 2206
rect 1898 2203 1908 2206
rect 1922 2203 1940 2206
rect 2042 2203 2068 2206
rect 2092 2203 2109 2206
rect 2122 2203 2132 2206
rect 2146 2203 2172 2206
rect 2514 2203 2532 2206
rect 2738 2203 2755 2206
rect 2844 2203 2861 2206
rect 3066 2203 3092 2206
rect 3122 2205 3125 2213
rect 3156 2203 3196 2206
rect 3236 2203 3261 2206
rect 3362 2203 3372 2206
rect 1058 2193 1076 2196
rect 1090 2193 1109 2196
rect 1434 2193 1444 2196
rect 1474 2193 1500 2196
rect 1546 2193 1564 2196
rect 1844 2193 1853 2196
rect 1962 2193 1972 2196
rect 2098 2193 2108 2196
rect 3138 2193 3148 2196
rect 38 2167 3434 2173
rect 380 2143 389 2146
rect 548 2143 565 2146
rect 1106 2143 1117 2146
rect 1218 2143 1244 2146
rect 1380 2143 1389 2146
rect 1474 2143 1492 2146
rect 1114 2136 1117 2143
rect 1618 2136 1621 2146
rect 1756 2143 1765 2146
rect 124 2133 133 2136
rect 194 2133 204 2136
rect 338 2133 364 2136
rect 482 2133 492 2136
rect 506 2133 532 2136
rect 546 2133 572 2136
rect 482 2126 485 2133
rect 618 2126 621 2134
rect 626 2133 652 2136
rect 690 2133 700 2136
rect 714 2133 756 2136
rect 810 2133 860 2136
rect 874 2133 884 2136
rect 908 2133 925 2136
rect 1042 2133 1076 2136
rect 1100 2133 1109 2136
rect 1114 2133 1124 2136
rect 1162 2133 1172 2136
rect 1204 2133 1252 2136
rect 1266 2133 1284 2136
rect 1308 2133 1333 2136
rect 1402 2133 1428 2136
rect 1452 2133 1461 2136
rect 1474 2133 1500 2136
rect 1538 2133 1588 2136
rect 1610 2133 1621 2136
rect 1716 2133 1733 2136
rect 1804 2133 1821 2136
rect 1842 2133 1845 2156
rect 2002 2153 2037 2156
rect 2002 2136 2005 2153
rect 2010 2143 2044 2146
rect 2146 2143 2156 2146
rect 2170 2143 2180 2146
rect 2274 2143 2300 2146
rect 2338 2143 2354 2146
rect 2482 2143 2500 2146
rect 2514 2143 2523 2146
rect 2636 2143 2645 2146
rect 1892 2133 1933 2136
rect 1954 2133 1972 2136
rect 1988 2133 2005 2136
rect 2026 2133 2051 2136
rect 2130 2133 2163 2136
rect 2188 2133 2205 2136
rect 2266 2133 2308 2136
rect 2364 2133 2381 2136
rect 98 2123 108 2126
rect 122 2123 133 2126
rect 130 2116 133 2123
rect 130 2113 164 2116
rect 170 2106 173 2125
rect 306 2123 324 2126
rect 346 2123 356 2126
rect 386 2123 404 2126
rect 474 2123 485 2126
rect 562 2123 580 2126
rect 618 2123 637 2126
rect 698 2123 708 2126
rect 714 2123 764 2126
rect 810 2123 852 2126
rect 876 2123 892 2126
rect 978 2123 997 2126
rect 978 2106 981 2123
rect 986 2113 1012 2116
rect 1036 2113 1069 2116
rect 1114 2106 1117 2133
rect 1122 2123 1132 2126
rect 1170 2123 1180 2126
rect 1260 2123 1269 2126
rect 146 2103 173 2106
rect 266 2103 284 2106
rect 978 2103 1028 2106
rect 1106 2103 1117 2106
rect 1266 2083 1269 2123
rect 1274 2123 1292 2126
rect 1338 2123 1356 2126
rect 1380 2123 1436 2126
rect 1524 2123 1533 2126
rect 1562 2123 1580 2126
rect 1610 2125 1613 2133
rect 1722 2123 1732 2126
rect 1756 2123 1765 2126
rect 1878 2123 1885 2126
rect 1930 2125 1933 2133
rect 2386 2126 2389 2134
rect 2402 2133 2420 2136
rect 2442 2133 2445 2143
rect 2466 2133 2501 2136
rect 2508 2133 2525 2136
rect 2532 2133 2565 2136
rect 2596 2133 2605 2136
rect 2634 2133 2676 2136
rect 2700 2133 2717 2136
rect 2722 2133 2732 2136
rect 2746 2127 2749 2136
rect 2874 2133 2884 2136
rect 3074 2133 3092 2136
rect 3164 2133 3181 2136
rect 3282 2133 3292 2136
rect 3356 2133 3364 2136
rect 1996 2123 2045 2126
rect 2076 2123 2085 2126
rect 2252 2123 2261 2126
rect 2316 2123 2325 2126
rect 2332 2123 2349 2126
rect 2378 2123 2389 2126
rect 2396 2123 2405 2126
rect 2460 2123 2477 2126
rect 2570 2123 2580 2126
rect 2636 2123 2645 2126
rect 2706 2123 2740 2126
rect 2746 2124 2764 2127
rect 2874 2126 2877 2133
rect 3282 2126 3285 2133
rect 2868 2123 2877 2126
rect 3004 2123 3029 2126
rect 3060 2123 3069 2126
rect 3220 2123 3229 2126
rect 3276 2123 3285 2126
rect 3362 2123 3372 2126
rect 1274 2113 1277 2123
rect 1308 2113 1317 2116
rect 1634 2113 1644 2116
rect 1716 2113 1725 2116
rect 1826 2113 1836 2116
rect 2082 2113 2091 2116
rect 2212 2113 2221 2116
rect 2756 2113 2765 2116
rect 2780 2113 2797 2116
rect 1626 2103 1660 2106
rect 1810 2103 1852 2106
rect 2210 2103 2228 2106
rect 14 2067 3458 2073
rect 3162 2053 3189 2056
rect 2578 2043 2613 2046
rect 162 2033 173 2036
rect 108 2023 133 2026
rect 170 2015 173 2033
rect 538 2023 549 2026
rect 546 2016 549 2023
rect 642 2016 645 2024
rect 650 2023 669 2026
rect 666 2016 669 2023
rect 194 2013 228 2016
rect 282 2013 332 2016
rect 372 2013 381 2016
rect 460 2013 469 2016
rect 474 2013 492 2016
rect 114 2003 140 2006
rect 218 2003 236 2006
rect 298 2003 324 2006
rect 410 2003 444 2006
rect 506 2005 509 2016
rect 516 2013 541 2016
rect 546 2013 564 2016
rect 602 2013 628 2016
rect 642 2013 661 2016
rect 666 2013 677 2016
rect 714 2013 748 2016
rect 786 2013 812 2016
rect 530 2003 556 2006
rect 580 2003 589 2006
rect 594 2003 620 2006
rect 644 2003 669 2006
rect 674 2005 677 2013
rect 708 2003 733 2006
rect 786 2003 804 2006
rect 850 1996 853 2036
rect 1482 2033 1493 2036
rect 2578 2033 2589 2036
rect 1314 2023 1349 2026
rect 1476 2023 1485 2026
rect 932 2013 941 2016
rect 946 2013 956 2016
rect 994 2013 1012 2016
rect 1034 2013 1076 2016
rect 1098 2013 1116 2016
rect 1138 2013 1148 2016
rect 1210 2013 1218 2016
rect 1244 2013 1261 2016
rect 1284 2013 1293 2016
rect 1308 2013 1341 2016
rect 1346 2006 1349 2023
rect 1370 2013 1380 2016
rect 858 2003 876 2006
rect 890 2003 908 2006
rect 1028 2003 1037 2006
rect 1042 2003 1068 2006
rect 1082 2003 1108 2006
rect 1122 2003 1140 2006
rect 1178 2003 1211 2006
rect 1226 2003 1236 2006
rect 1242 2003 1276 2006
rect 1306 2003 1349 2006
rect 1354 2003 1372 2006
rect 1442 2003 1452 2006
rect 372 1993 389 1996
rect 850 1993 868 1996
rect 962 1993 997 1996
rect 1490 1986 1493 2033
rect 1836 2023 1853 2026
rect 1884 2023 1909 2026
rect 2188 2023 2205 2026
rect 1674 2013 1725 2016
rect 1780 2013 1789 2016
rect 1794 2013 1820 2016
rect 1882 2013 1932 2016
rect 1988 2013 1997 2016
rect 2010 2013 2020 2016
rect 2052 2013 2077 2016
rect 2162 2013 2172 2016
rect 2284 2013 2309 2016
rect 2316 2013 2333 2016
rect 1674 2006 1677 2013
rect 1498 2003 1532 2006
rect 1564 2003 1581 2006
rect 1594 2003 1620 2006
rect 1642 2003 1660 2006
rect 1666 2003 1677 2006
rect 1722 2003 1725 2013
rect 1740 2003 1756 2006
rect 1786 1996 1789 2013
rect 1836 2003 1845 2006
rect 1882 2005 1885 2013
rect 1954 2003 1980 2006
rect 2058 2003 2100 2006
rect 2132 2003 2163 2006
rect 2188 2003 2197 2006
rect 2202 2003 2228 2006
rect 2276 2003 2293 2006
rect 2298 2003 2308 2006
rect 2380 2003 2397 2006
rect 2412 2003 2445 2006
rect 2452 2003 2469 2006
rect 2476 2003 2509 2006
rect 1786 1993 1797 1996
rect 1954 1993 1972 1996
rect 2210 1993 2220 1996
rect 2322 1993 2348 1996
rect 2418 1993 2444 1996
rect 2458 1993 2468 1996
rect 650 1983 669 1986
rect 1490 1983 1525 1986
rect 2514 1983 2517 2026
rect 2586 2016 2589 2033
rect 2522 2013 2532 2016
rect 2578 2013 2589 2016
rect 2594 2013 2628 2016
rect 2578 2006 2581 2013
rect 2658 2006 2661 2036
rect 2778 2013 2795 2016
rect 2826 2013 2852 2016
rect 2890 2013 2908 2016
rect 2932 2013 2941 2016
rect 2954 2013 2964 2016
rect 3028 2013 3061 2016
rect 3106 2013 3132 2016
rect 3292 2013 3317 2016
rect 2572 2003 2581 2006
rect 2586 2003 2620 2006
rect 2658 2003 2676 2006
rect 2730 2003 2740 2006
rect 2756 2003 2765 2006
rect 2818 2003 2843 2006
rect 2906 2003 2916 2006
rect 2930 2003 2956 2006
rect 2970 2003 3012 2006
rect 3026 2003 3060 2006
rect 3098 2003 3140 2006
rect 2586 1996 2589 2003
rect 2578 1993 2589 1996
rect 2932 1993 2941 1996
rect 3028 1993 3053 1996
rect 38 1967 3434 1973
rect 124 1923 133 1926
rect 162 1923 180 1926
rect 186 1923 196 1926
rect 218 1916 221 1936
rect 234 1925 237 1956
rect 1018 1953 1045 1956
rect 692 1943 709 1946
rect 946 1943 957 1946
rect 1066 1943 1084 1946
rect 514 1926 517 1936
rect 554 1926 557 1934
rect 562 1933 572 1936
rect 642 1933 676 1936
rect 746 1933 788 1936
rect 810 1933 828 1936
rect 842 1933 876 1936
rect 932 1933 949 1936
rect 954 1926 957 1943
rect 1234 1936 1237 1945
rect 1330 1936 1333 1956
rect 1514 1943 1556 1946
rect 1794 1936 1797 1956
rect 1834 1953 1845 1956
rect 1842 1936 1845 1953
rect 1938 1943 1972 1946
rect 2082 1943 2091 1946
rect 962 1933 972 1936
rect 1004 1933 1045 1936
rect 1092 1933 1117 1936
rect 1178 1933 1196 1936
rect 1228 1933 1237 1936
rect 1250 1933 1284 1936
rect 1308 1933 1333 1936
rect 1386 1933 1396 1936
rect 1514 1933 1581 1936
rect 1620 1933 1645 1936
rect 1658 1933 1668 1936
rect 1794 1933 1804 1936
rect 1842 1933 1859 1936
rect 1890 1933 1901 1936
rect 1924 1933 1957 1936
rect 2090 1933 2100 1936
rect 2106 1933 2115 1936
rect 2156 1933 2181 1936
rect 290 1923 308 1926
rect 314 1923 324 1926
rect 396 1923 405 1926
rect 412 1923 437 1926
rect 514 1923 540 1926
rect 554 1923 573 1926
rect 580 1923 597 1926
rect 602 1923 620 1926
rect 810 1923 836 1926
rect 890 1923 916 1926
rect 954 1923 980 1926
rect 1026 1923 1060 1926
rect 108 1913 117 1916
rect 132 1913 165 1916
rect 204 1913 221 1916
rect 252 1913 261 1916
rect 340 1913 349 1916
rect 402 1913 405 1923
rect 468 1913 477 1916
rect 508 1913 517 1916
rect 556 1913 565 1916
rect 636 1913 661 1916
rect 932 1913 941 1916
rect 1114 1906 1117 1933
rect 1890 1926 1893 1933
rect 1186 1923 1204 1926
rect 1274 1923 1292 1926
rect 1306 1923 1348 1926
rect 1394 1923 1404 1926
rect 1508 1923 1533 1926
rect 1572 1923 1589 1926
rect 1676 1923 1685 1926
rect 1834 1923 1867 1926
rect 1882 1923 1893 1926
rect 1932 1923 1973 1926
rect 1994 1923 2004 1926
rect 1882 1916 1885 1923
rect 2090 1922 2093 1933
rect 2194 1926 2197 1943
rect 2210 1936 2213 1946
rect 2666 1943 2683 1946
rect 3124 1943 3133 1946
rect 2204 1933 2213 1936
rect 2316 1933 2341 1936
rect 2388 1933 2397 1936
rect 2404 1933 2437 1936
rect 2442 1926 2445 1934
rect 2498 1926 2501 1934
rect 2164 1923 2197 1926
rect 2266 1923 2284 1926
rect 2418 1923 2445 1926
rect 2490 1923 2501 1926
rect 2530 1925 2533 1936
rect 2554 1933 2564 1936
rect 2590 1933 2613 1936
rect 2650 1933 2660 1936
rect 2666 1933 2692 1936
rect 2698 1933 2732 1936
rect 2788 1933 2821 1936
rect 2490 1916 2493 1923
rect 1132 1913 1141 1916
rect 1364 1913 1389 1916
rect 1828 1913 1837 1916
rect 2052 1913 2085 1916
rect 2482 1913 2493 1916
rect 2514 1913 2523 1916
rect 2610 1906 2613 1933
rect 2826 1926 2829 1934
rect 2876 1933 2917 1936
rect 2922 1926 2925 1934
rect 2938 1933 2948 1936
rect 2954 1933 2964 1936
rect 3012 1933 3037 1936
rect 3060 1933 3085 1936
rect 2668 1923 2685 1926
rect 2722 1923 2740 1926
rect 2786 1923 2829 1926
rect 2890 1923 2925 1926
rect 3020 1923 3029 1926
rect 3034 1925 3037 1933
rect 3124 1923 3133 1926
rect 3244 1923 3269 1926
rect 3396 1923 3469 1926
rect 2620 1913 2629 1916
rect 218 1903 244 1906
rect 426 1903 460 1906
rect 1114 1903 1148 1906
rect 2530 1903 2539 1906
rect 2610 1903 2621 1906
rect 14 1867 3458 1873
rect 3466 1856 3469 1923
rect 3370 1853 3469 1856
rect 250 1833 261 1836
rect 378 1833 397 1836
rect 196 1823 205 1826
rect 82 1813 100 1816
rect 170 1813 180 1816
rect 258 1815 261 1833
rect 332 1823 341 1826
rect 356 1823 365 1826
rect 394 1815 397 1833
rect 458 1813 484 1816
rect 132 1803 165 1806
rect 458 1803 461 1813
rect 490 1806 493 1825
rect 530 1816 533 1825
rect 756 1823 789 1826
rect 820 1823 829 1826
rect 868 1823 877 1826
rect 956 1823 989 1826
rect 1036 1823 1077 1826
rect 1108 1823 1157 1826
rect 1444 1823 1469 1826
rect 1692 1823 1725 1826
rect 2298 1823 2317 1826
rect 2484 1823 2517 1826
rect 2538 1825 2541 1836
rect 2626 1833 2645 1836
rect 2698 1833 2755 1836
rect 2914 1833 2924 1836
rect 2596 1823 2605 1826
rect 2610 1823 2636 1826
rect 1722 1816 1725 1823
rect 2642 1816 2645 1833
rect 2692 1823 2701 1826
rect 2802 1823 2813 1826
rect 2932 1823 2941 1826
rect 3020 1823 3029 1826
rect 498 1813 524 1816
rect 530 1813 541 1816
rect 572 1813 581 1816
rect 668 1813 677 1816
rect 770 1813 804 1816
rect 826 1813 860 1816
rect 994 1813 1020 1816
rect 1082 1813 1092 1816
rect 1228 1813 1237 1816
rect 1338 1813 1356 1816
rect 1442 1813 1453 1816
rect 1514 1813 1549 1816
rect 1722 1813 1733 1816
rect 1740 1813 1749 1816
rect 1818 1813 1836 1816
rect 1954 1813 1972 1816
rect 2052 1813 2061 1816
rect 2092 1813 2101 1816
rect 2106 1813 2132 1816
rect 2154 1813 2172 1816
rect 2258 1813 2268 1816
rect 2298 1813 2340 1816
rect 2354 1813 2372 1816
rect 2386 1813 2429 1816
rect 466 1803 476 1806
rect 490 1803 501 1806
rect 634 1803 660 1806
rect 778 1803 796 1806
rect 866 1803 908 1806
rect 956 1803 997 1806
rect 1050 1803 1084 1806
rect 1122 1803 1156 1806
rect 1186 1803 1204 1806
rect 1242 1803 1276 1806
rect 1300 1803 1341 1806
rect 498 1793 501 1803
rect 1450 1796 1453 1813
rect 1500 1803 1541 1806
rect 1546 1805 1549 1813
rect 1572 1803 1629 1806
rect 1650 1803 1676 1806
rect 1698 1803 1732 1806
rect 1756 1803 1789 1806
rect 1818 1803 1828 1806
rect 1866 1803 1916 1806
rect 1978 1803 2012 1806
rect 2036 1803 2044 1806
rect 2114 1803 2124 1806
rect 2188 1803 2197 1806
rect 2306 1803 2332 1806
rect 2388 1803 2421 1806
rect 2426 1805 2429 1813
rect 2450 1813 2461 1816
rect 2796 1813 2805 1816
rect 2810 1813 2813 1823
rect 3250 1816 3253 1826
rect 3332 1823 3341 1826
rect 3338 1816 3341 1823
rect 2858 1813 2876 1816
rect 2954 1813 2972 1816
rect 2994 1813 3003 1816
rect 3034 1813 3092 1816
rect 3138 1813 3164 1816
rect 3170 1813 3196 1816
rect 3236 1813 3253 1816
rect 3314 1813 3323 1816
rect 3338 1813 3356 1816
rect 2450 1805 2453 1813
rect 2484 1803 2509 1806
rect 2692 1803 2725 1806
rect 1450 1793 1492 1796
rect 1586 1793 1628 1796
rect 2194 1793 2213 1796
rect 2746 1783 2749 1813
rect 2818 1803 2835 1806
rect 2914 1803 2917 1813
rect 3034 1803 3037 1813
rect 3130 1803 3156 1806
rect 3170 1803 3173 1813
rect 3202 1803 3220 1806
rect 3250 1803 3292 1806
rect 38 1767 3434 1773
rect 906 1743 933 1746
rect 1634 1743 1660 1746
rect 1954 1743 1964 1746
rect 2162 1743 2189 1746
rect 3106 1743 3117 1746
rect 66 1733 84 1736
rect 162 1733 172 1736
rect 194 1733 220 1736
rect 242 1733 252 1736
rect 282 1733 300 1736
rect 354 1726 357 1734
rect 386 1733 404 1736
rect 522 1733 532 1736
rect 594 1733 636 1736
rect 700 1733 717 1736
rect 730 1733 740 1736
rect 890 1733 948 1736
rect 1154 1733 1196 1736
rect 1258 1733 1284 1736
rect 106 1723 124 1726
rect 154 1723 164 1726
rect 202 1723 212 1726
rect 298 1723 308 1726
rect 354 1723 373 1726
rect 378 1723 412 1726
rect 444 1723 453 1726
rect 522 1723 525 1733
rect 1306 1726 1309 1734
rect 1314 1733 1372 1736
rect 1396 1733 1413 1736
rect 1418 1733 1436 1736
rect 1450 1733 1500 1736
rect 1514 1733 1532 1736
rect 1546 1733 1596 1736
rect 1650 1733 1668 1736
rect 1722 1733 1732 1736
rect 610 1723 643 1726
rect 666 1723 684 1726
rect 132 1713 149 1716
rect 154 1693 157 1723
rect 370 1716 373 1723
rect 356 1713 365 1716
rect 370 1713 381 1716
rect 564 1713 573 1716
rect 588 1713 637 1716
rect 666 1713 669 1723
rect 802 1713 812 1716
rect 818 1706 821 1725
rect 842 1723 884 1726
rect 972 1723 989 1726
rect 1178 1723 1204 1726
rect 1306 1723 1373 1726
rect 1394 1723 1444 1726
rect 1466 1723 1508 1726
rect 1530 1723 1540 1726
rect 1554 1723 1604 1726
rect 1650 1716 1653 1733
rect 1754 1726 1757 1734
rect 1850 1733 1860 1736
rect 1898 1733 1916 1736
rect 1940 1733 1965 1736
rect 2050 1733 2060 1736
rect 2122 1733 2132 1736
rect 2162 1726 2165 1743
rect 3106 1736 3109 1743
rect 2170 1734 2196 1736
rect 2170 1733 2197 1734
rect 2210 1733 2228 1736
rect 1676 1723 1685 1726
rect 1706 1723 1740 1726
rect 1754 1723 1773 1726
rect 1884 1723 1901 1726
rect 1914 1723 1924 1726
rect 1988 1723 1997 1726
rect 2010 1723 2028 1726
rect 2076 1723 2093 1726
rect 2106 1723 2115 1726
rect 2162 1723 2173 1726
rect 2194 1723 2197 1733
rect 2266 1726 2269 1734
rect 2388 1733 2405 1736
rect 2476 1733 2493 1736
rect 2540 1733 2557 1736
rect 2590 1733 2613 1736
rect 2684 1733 2701 1736
rect 2764 1733 2781 1736
rect 2804 1733 2821 1736
rect 2826 1733 2853 1736
rect 2204 1723 2229 1726
rect 2250 1723 2269 1726
rect 2290 1723 2340 1726
rect 2354 1723 2372 1726
rect 2394 1723 2428 1726
rect 2596 1723 2637 1726
rect 836 1713 853 1716
rect 892 1713 917 1716
rect 1028 1713 1037 1716
rect 1052 1713 1061 1716
rect 1124 1713 1133 1716
rect 1148 1713 1189 1716
rect 1220 1713 1237 1716
rect 1396 1713 1405 1716
rect 1452 1713 1493 1716
rect 1620 1713 1653 1716
rect 1756 1713 1765 1716
rect 1770 1706 1773 1723
rect 2698 1716 2701 1733
rect 2850 1726 2853 1733
rect 2930 1733 2941 1736
rect 2954 1733 2964 1736
rect 2980 1733 3013 1736
rect 3100 1733 3109 1736
rect 3114 1733 3140 1736
rect 3194 1733 3228 1736
rect 2930 1726 2933 1733
rect 3378 1726 3381 1734
rect 2706 1723 2747 1726
rect 2762 1723 2780 1726
rect 2812 1723 2845 1726
rect 2850 1723 2868 1726
rect 2924 1723 2933 1726
rect 2988 1723 3021 1726
rect 3074 1723 3084 1726
rect 3130 1723 3148 1726
rect 3268 1723 3293 1726
rect 3330 1723 3364 1726
rect 3378 1723 3405 1726
rect 1786 1713 1804 1716
rect 1828 1713 1837 1716
rect 2292 1713 2325 1716
rect 2698 1713 2709 1716
rect 562 1703 580 1706
rect 762 1703 821 1706
rect 994 1703 1044 1706
rect 1770 1703 1820 1706
rect 2322 1703 2325 1713
rect 3290 1706 3293 1723
rect 3324 1713 3349 1716
rect 3380 1713 3397 1716
rect 3402 1706 3405 1723
rect 3290 1703 3316 1706
rect 3394 1703 3405 1706
rect 594 1683 629 1686
rect 2818 1683 2853 1686
rect 14 1667 3458 1673
rect 578 1633 597 1636
rect 1146 1633 1165 1636
rect 1626 1633 1653 1636
rect 1890 1633 1893 1656
rect 2858 1643 2885 1646
rect 3370 1643 3397 1646
rect 148 1623 181 1626
rect 562 1623 588 1626
rect 122 1613 133 1616
rect 140 1613 149 1616
rect 170 1613 188 1616
rect 282 1613 292 1616
rect 324 1615 333 1616
rect 322 1613 333 1615
rect 420 1613 468 1616
rect 482 1613 501 1616
rect 556 1613 565 1616
rect 594 1615 597 1633
rect 612 1623 629 1626
rect 780 1623 813 1626
rect 1122 1623 1156 1626
rect 626 1613 652 1616
rect 746 1613 764 1616
rect 778 1613 836 1616
rect 892 1613 901 1616
rect 906 1613 940 1616
rect 972 1613 989 1616
rect 994 1613 1028 1616
rect 1052 1613 1093 1616
rect 1100 1613 1141 1616
rect 1162 1615 1165 1633
rect 1180 1623 1197 1626
rect 1500 1623 1509 1626
rect 1620 1623 1645 1626
rect 1218 1613 1228 1616
rect 1314 1613 1332 1616
rect 1346 1613 1396 1616
rect 130 1606 133 1613
rect 322 1606 325 1613
rect 482 1606 485 1613
rect 1642 1606 1645 1623
rect 1650 1616 1653 1633
rect 1796 1623 1805 1626
rect 1890 1623 1909 1626
rect 1980 1623 1997 1626
rect 1890 1616 1893 1623
rect 2122 1616 2125 1636
rect 2396 1623 2413 1626
rect 2460 1623 2477 1626
rect 2508 1623 2541 1626
rect 2818 1616 2821 1636
rect 3298 1633 3325 1636
rect 3082 1623 3093 1626
rect 3274 1623 3316 1626
rect 1650 1613 1660 1616
rect 1706 1613 1740 1616
rect 1842 1613 1852 1616
rect 1884 1613 1893 1616
rect 1898 1613 1916 1616
rect 1954 1613 1964 1616
rect 2010 1613 2036 1616
rect 2050 1613 2061 1616
rect 2066 1613 2084 1616
rect 2122 1613 2133 1616
rect 2188 1613 2205 1616
rect 2220 1613 2229 1616
rect 2242 1613 2252 1616
rect 2340 1613 2373 1616
rect 2394 1613 2444 1616
rect 2458 1613 2485 1616
rect 2530 1613 2548 1616
rect 2580 1613 2597 1616
rect 2666 1613 2684 1616
rect 2698 1613 2716 1616
rect 2730 1613 2757 1616
rect 2770 1613 2780 1616
rect 2818 1613 2829 1616
rect 2890 1613 2900 1616
rect 3004 1613 3021 1616
rect 3060 1613 3085 1616
rect 74 1603 100 1606
rect 212 1603 221 1606
rect 226 1603 236 1606
rect 258 1603 293 1606
rect 322 1603 356 1606
rect 372 1603 381 1606
rect 386 1603 412 1606
rect 434 1603 460 1606
rect 498 1603 532 1606
rect 708 1603 741 1606
rect 858 1603 884 1606
rect 938 1603 948 1606
rect 964 1603 973 1606
rect 986 1603 1036 1606
rect 1050 1603 1092 1606
rect 1202 1603 1236 1606
rect 1306 1603 1324 1606
rect 1348 1603 1373 1606
rect 1378 1603 1404 1606
rect 1420 1603 1437 1606
rect 1442 1603 1476 1606
rect 1500 1603 1525 1606
rect 1564 1603 1581 1606
rect 1642 1603 1668 1606
rect 1722 1603 1732 1606
rect 1802 1603 1859 1606
rect 1882 1603 1908 1606
rect 1986 1603 1996 1606
rect 2050 1605 2053 1613
rect 74 1583 77 1603
rect 2066 1593 2069 1613
rect 2130 1606 2133 1613
rect 2074 1603 2091 1606
rect 2194 1603 2212 1606
rect 2276 1603 2285 1606
rect 2290 1603 2316 1606
rect 2346 1603 2372 1606
rect 2458 1605 2461 1613
rect 2754 1606 2757 1613
rect 2826 1606 2829 1613
rect 2466 1603 2484 1606
rect 2514 1603 2556 1606
rect 2572 1603 2581 1606
rect 2628 1603 2637 1606
rect 2650 1603 2676 1606
rect 2700 1603 2708 1606
rect 2732 1603 2749 1606
rect 2754 1603 2788 1606
rect 2852 1603 2892 1606
rect 2956 1603 2989 1606
rect 3010 1603 3036 1606
rect 3042 1603 3052 1606
rect 3090 1603 3093 1623
rect 3322 1616 3325 1633
rect 3364 1623 3397 1626
rect 3172 1613 3181 1616
rect 3234 1603 3244 1606
rect 2074 1586 2077 1603
rect 3210 1593 3220 1596
rect 2058 1583 2077 1586
rect 2642 1583 2661 1586
rect 38 1567 3434 1573
rect 330 1536 333 1556
rect 1426 1553 1469 1556
rect 1866 1553 1893 1556
rect 3034 1546 3037 1556
rect 498 1536 501 1546
rect 106 1533 116 1536
rect 130 1533 148 1536
rect 164 1533 173 1536
rect 236 1533 245 1536
rect 330 1533 362 1536
rect 380 1533 389 1536
rect 450 1533 460 1536
rect 498 1533 532 1536
rect 642 1533 660 1536
rect 690 1533 708 1536
rect 788 1533 805 1536
rect 858 1533 868 1536
rect 884 1533 893 1536
rect 130 1526 133 1533
rect 498 1526 501 1533
rect 930 1526 933 1534
rect 986 1533 997 1536
rect 1020 1533 1077 1536
rect 1172 1533 1181 1536
rect 1186 1533 1236 1536
rect 1258 1533 1308 1536
rect 1346 1533 1372 1536
rect 1420 1533 1453 1536
rect 986 1526 989 1533
rect 1474 1526 1477 1546
rect 1738 1536 1741 1546
rect 2210 1543 2221 1546
rect 2218 1536 2221 1543
rect 2458 1543 2477 1546
rect 3034 1543 3060 1546
rect 2458 1536 2461 1543
rect 1738 1533 1755 1536
rect 1794 1533 1804 1536
rect 1924 1533 1933 1536
rect 82 1523 100 1526
rect 124 1523 133 1526
rect 178 1523 212 1526
rect 250 1523 260 1526
rect 274 1523 292 1526
rect 330 1523 355 1526
rect 418 1523 444 1526
rect 468 1523 501 1526
rect 556 1523 581 1526
rect 684 1523 709 1526
rect 718 1523 757 1526
rect 842 1523 860 1526
rect 898 1523 933 1526
rect 940 1523 989 1526
rect 1028 1523 1037 1526
rect 1138 1523 1156 1526
rect 1260 1523 1285 1526
rect 1380 1523 1404 1526
rect 1474 1523 1492 1526
rect 1546 1523 1556 1526
rect 1570 1523 1620 1526
rect 1738 1523 1764 1526
rect 1786 1523 1812 1526
rect 1818 1523 1828 1526
rect 418 1513 421 1523
rect 476 1513 517 1516
rect 628 1513 653 1516
rect 1084 1513 1093 1516
rect 1108 1513 1125 1516
rect 1572 1513 1581 1516
rect 1666 1513 1700 1516
rect 1938 1513 1941 1534
rect 1954 1533 1989 1536
rect 2020 1533 2029 1536
rect 2066 1533 2091 1536
rect 2146 1533 2180 1536
rect 2196 1533 2213 1536
rect 2218 1533 2236 1536
rect 2394 1533 2420 1536
rect 2436 1533 2461 1536
rect 2466 1533 2492 1536
rect 2508 1533 2517 1536
rect 2562 1533 2580 1536
rect 2668 1533 2708 1536
rect 2730 1533 2805 1536
rect 2812 1533 2845 1536
rect 2884 1533 2893 1536
rect 2906 1533 2916 1536
rect 2954 1533 2973 1536
rect 3028 1533 3037 1536
rect 3042 1533 3061 1536
rect 3106 1533 3116 1536
rect 1986 1526 1989 1533
rect 1948 1523 1981 1526
rect 1986 1523 1996 1526
rect 2034 1523 2044 1526
rect 2066 1516 2069 1533
rect 2074 1523 2100 1526
rect 2132 1523 2141 1526
rect 2260 1523 2301 1526
rect 2330 1523 2340 1526
rect 2516 1523 2525 1526
rect 2538 1523 2572 1526
rect 2690 1523 2700 1526
rect 2730 1525 2733 1533
rect 3138 1526 3141 1534
rect 3290 1533 3323 1536
rect 3346 1533 3356 1536
rect 3394 1533 3405 1536
rect 2796 1523 2805 1526
rect 2882 1523 2924 1526
rect 2970 1523 2980 1526
rect 3084 1523 3093 1526
rect 3124 1523 3141 1526
rect 3306 1523 3332 1526
rect 3346 1523 3364 1526
rect 1956 1513 1965 1516
rect 2052 1513 2061 1516
rect 2066 1513 2077 1516
rect 1658 1503 1716 1506
rect 2138 1493 2141 1523
rect 2356 1513 2365 1516
rect 2884 1513 2893 1516
rect 3156 1513 3165 1516
rect 3228 1513 3253 1516
rect 3258 1506 3261 1515
rect 3284 1513 3325 1516
rect 3373 1513 3397 1516
rect 3194 1503 3220 1506
rect 3234 1503 3261 1506
rect 3378 1503 3397 1506
rect 3402 1496 3405 1533
rect 3378 1493 3405 1496
rect 826 1483 853 1486
rect 946 1483 989 1486
rect 14 1467 3458 1473
rect 244 1423 253 1426
rect 82 1413 100 1416
rect 226 1413 236 1416
rect 116 1403 125 1406
rect 130 1403 140 1406
rect 164 1403 181 1406
rect 130 1396 133 1403
rect 122 1393 133 1396
rect 274 1386 277 1436
rect 330 1416 333 1446
rect 330 1413 340 1416
rect 378 1406 381 1426
rect 386 1416 389 1446
rect 482 1416 485 1456
rect 666 1443 677 1446
rect 722 1443 749 1446
rect 386 1413 411 1416
rect 460 1413 477 1416
rect 482 1413 500 1416
rect 426 1406 429 1413
rect 474 1406 477 1413
rect 282 1403 300 1406
rect 316 1403 333 1406
rect 378 1403 404 1406
rect 418 1403 429 1406
rect 452 1403 469 1406
rect 474 1403 508 1406
rect 274 1383 285 1386
rect 330 1383 333 1403
rect 466 1396 469 1403
rect 466 1393 485 1396
rect 538 1383 541 1436
rect 562 1433 572 1436
rect 594 1433 613 1436
rect 546 1423 556 1426
rect 594 1396 597 1433
rect 602 1413 620 1416
rect 666 1406 669 1443
rect 722 1416 725 1443
rect 930 1433 964 1436
rect 2994 1433 3020 1436
rect 718 1413 725 1416
rect 730 1413 756 1416
rect 794 1406 797 1426
rect 930 1423 948 1426
rect 972 1423 981 1426
rect 1036 1423 1061 1426
rect 1100 1423 1125 1426
rect 1460 1423 1485 1426
rect 1652 1423 1685 1426
rect 1804 1423 1853 1426
rect 2228 1423 2245 1426
rect 2860 1423 2869 1426
rect 836 1413 900 1416
rect 1028 1413 1084 1416
rect 1098 1413 1156 1416
rect 1266 1413 1325 1416
rect 1380 1413 1389 1416
rect 1410 1413 1444 1416
rect 1530 1413 1572 1416
rect 1610 1413 1644 1416
rect 1690 1413 1700 1416
rect 1810 1413 1868 1416
rect 1940 1413 1957 1416
rect 1964 1413 1981 1416
rect 2178 1413 2212 1416
rect 2226 1413 2268 1416
rect 2322 1413 2348 1416
rect 2370 1413 2404 1416
rect 2514 1413 2532 1416
rect 2602 1413 2612 1416
rect 2658 1413 2676 1416
rect 2706 1413 2717 1416
rect 2796 1413 2837 1416
rect 2964 1413 2973 1416
rect 1322 1406 1325 1413
rect 2706 1406 2709 1413
rect 2994 1406 2997 1433
rect 3028 1423 3045 1426
rect 3124 1423 3133 1426
rect 3244 1423 3253 1426
rect 3316 1423 3325 1426
rect 3034 1413 3052 1416
rect 3082 1413 3108 1416
rect 3180 1413 3205 1416
rect 3282 1413 3300 1416
rect 3338 1413 3364 1416
rect 610 1403 628 1406
rect 644 1403 669 1406
rect 708 1403 733 1406
rect 780 1403 797 1406
rect 802 1403 828 1406
rect 858 1403 892 1406
rect 916 1403 925 1406
rect 1010 1403 1020 1406
rect 1100 1403 1117 1406
rect 1122 1403 1164 1406
rect 1274 1403 1284 1406
rect 1322 1403 1356 1406
rect 1372 1403 1381 1406
rect 1426 1403 1436 1406
rect 1460 1403 1485 1406
rect 1500 1403 1525 1406
rect 1546 1403 1564 1406
rect 1658 1403 1692 1406
rect 1804 1403 1853 1406
rect 1884 1403 1909 1406
rect 1946 1403 1956 1406
rect 1970 1403 2004 1406
rect 2100 1403 2140 1406
rect 2378 1403 2396 1406
rect 2436 1403 2453 1406
rect 2466 1403 2492 1406
rect 2498 1403 2524 1406
rect 2538 1403 2604 1406
rect 2650 1403 2668 1406
rect 2692 1403 2709 1406
rect 2746 1403 2788 1406
rect 2810 1403 2836 1406
rect 2860 1403 2901 1406
rect 2956 1403 2997 1406
rect 3074 1403 3100 1406
rect 3154 1403 3172 1406
rect 3186 1403 3220 1406
rect 3244 1403 3253 1406
rect 3258 1403 3292 1406
rect 3316 1403 3341 1406
rect 594 1393 613 1396
rect 2066 1393 2092 1396
rect 2410 1393 2428 1396
rect 2458 1393 2484 1396
rect 2538 1393 2541 1403
rect 2882 1393 2900 1396
rect 2930 1393 2948 1396
rect 3346 1383 3349 1413
rect 38 1367 3434 1373
rect 362 1343 381 1346
rect 546 1336 549 1356
rect 786 1353 805 1356
rect 802 1336 805 1353
rect 850 1343 861 1346
rect 978 1343 997 1346
rect 1330 1343 1341 1346
rect 82 1333 92 1336
rect 210 1333 236 1336
rect 260 1333 293 1336
rect 316 1333 333 1336
rect 538 1333 549 1336
rect 698 1333 724 1336
rect 772 1333 781 1336
rect 802 1333 811 1336
rect 836 1333 853 1336
rect 90 1323 100 1326
rect 138 1323 148 1326
rect 180 1323 221 1326
rect 226 1323 244 1326
rect 324 1323 333 1326
rect 396 1323 420 1326
rect 514 1323 532 1326
rect 636 1323 653 1326
rect 108 1313 125 1316
rect 138 1303 141 1323
rect 698 1316 701 1333
rect 732 1323 756 1326
rect 810 1323 820 1326
rect 260 1313 285 1316
rect 436 1313 445 1316
rect 540 1313 565 1316
rect 660 1313 669 1316
rect 684 1313 701 1316
rect 772 1313 797 1316
rect 562 1283 565 1313
rect 690 1303 709 1306
rect 690 1293 693 1303
rect 858 1286 861 1343
rect 1338 1336 1341 1343
rect 1858 1343 1877 1346
rect 2244 1343 2253 1346
rect 2354 1343 2372 1346
rect 2554 1343 2572 1346
rect 892 1333 901 1336
rect 914 1333 932 1336
rect 956 1333 965 1336
rect 978 1333 1004 1336
rect 1028 1333 1061 1336
rect 1092 1333 1101 1336
rect 1130 1333 1140 1336
rect 1244 1333 1261 1336
rect 1266 1333 1300 1336
rect 1324 1333 1333 1336
rect 1338 1333 1381 1336
rect 1388 1333 1429 1336
rect 906 1323 940 1326
rect 954 1323 973 1326
rect 954 1315 957 1323
rect 1028 1313 1045 1316
rect 1058 1313 1061 1333
rect 1266 1326 1269 1333
rect 1434 1326 1437 1335
rect 1546 1333 1596 1336
rect 1620 1333 1637 1336
rect 1682 1333 1741 1336
rect 1764 1333 1805 1336
rect 1810 1333 1820 1336
rect 1802 1326 1805 1333
rect 1858 1326 1861 1343
rect 3282 1336 3285 1346
rect 3394 1336 3397 1356
rect 1908 1333 1941 1336
rect 1946 1326 1949 1335
rect 1114 1323 1148 1326
rect 1250 1323 1269 1326
rect 1274 1323 1308 1326
rect 1396 1323 1405 1326
rect 1410 1323 1437 1326
rect 1444 1323 1477 1326
rect 1482 1323 1516 1326
rect 1546 1323 1604 1326
rect 1730 1323 1740 1326
rect 1772 1323 1789 1326
rect 1802 1323 1861 1326
rect 1874 1323 1884 1326
rect 1916 1323 1925 1326
rect 1930 1323 1949 1326
rect 2026 1326 2029 1335
rect 2034 1333 2068 1336
rect 2146 1333 2156 1336
rect 2380 1333 2405 1336
rect 2452 1333 2500 1336
rect 2532 1333 2596 1336
rect 2610 1333 2644 1336
rect 2674 1333 2692 1336
rect 2730 1333 2740 1336
rect 2764 1333 2773 1336
rect 2778 1333 2804 1336
rect 2828 1333 2853 1336
rect 2892 1333 2909 1336
rect 2954 1333 2988 1336
rect 3130 1333 3140 1336
rect 3170 1333 3204 1336
rect 3234 1333 3244 1336
rect 3282 1333 3300 1336
rect 3324 1333 3333 1336
rect 3346 1333 3356 1336
rect 3380 1333 3397 1336
rect 2906 1326 2909 1333
rect 3282 1326 3285 1333
rect 2026 1323 2037 1326
rect 2042 1323 2060 1326
rect 2098 1323 2148 1326
rect 2202 1323 2220 1326
rect 2274 1323 2292 1326
rect 2298 1323 2340 1326
rect 2388 1323 2397 1326
rect 2418 1323 2428 1326
rect 2458 1323 2508 1326
rect 2652 1323 2661 1326
rect 2682 1323 2700 1326
rect 2906 1323 2924 1326
rect 2938 1323 2996 1326
rect 3114 1323 3148 1326
rect 3202 1323 3212 1326
rect 3252 1323 3285 1326
rect 3354 1323 3364 1326
rect 1474 1316 1477 1323
rect 1092 1313 1125 1316
rect 1474 1313 1485 1316
rect 1532 1313 1589 1316
rect 1620 1313 1645 1316
rect 1676 1313 1725 1316
rect 1730 1306 1733 1323
rect 2660 1313 2677 1316
rect 2716 1313 2733 1316
rect 2764 1313 2773 1316
rect 3028 1313 3037 1316
rect 3042 1313 3084 1316
rect 3108 1313 3133 1316
rect 3164 1313 3173 1316
rect 3220 1313 3229 1316
rect 3260 1313 3277 1316
rect 1722 1303 1733 1306
rect 3034 1306 3037 1313
rect 3034 1303 3061 1306
rect 850 1283 861 1286
rect 14 1267 3458 1273
rect 1298 1253 1317 1256
rect 242 1243 253 1246
rect 170 1216 173 1236
rect 250 1223 253 1243
rect 322 1216 325 1236
rect 442 1226 445 1246
rect 1018 1243 1061 1246
rect 372 1223 405 1226
rect 420 1223 445 1226
rect 476 1223 509 1226
rect 644 1223 653 1226
rect 764 1223 781 1226
rect 828 1223 837 1226
rect 908 1223 949 1226
rect 506 1216 509 1223
rect 74 1213 100 1216
rect 156 1213 165 1216
rect 170 1213 204 1216
rect 250 1213 284 1216
rect 322 1213 362 1216
rect 378 1213 411 1216
rect 450 1213 460 1216
rect 506 1213 517 1216
rect 538 1213 588 1216
rect 602 1213 635 1216
rect 650 1213 653 1223
rect 658 1213 692 1216
rect 778 1213 781 1223
rect 794 1213 805 1216
rect 834 1213 853 1216
rect 946 1213 980 1216
rect 74 1203 77 1213
rect 658 1206 661 1213
rect 802 1206 805 1213
rect 1050 1206 1053 1236
rect 1058 1216 1061 1243
rect 1498 1233 1556 1236
rect 1746 1233 1756 1236
rect 1778 1233 1829 1236
rect 1906 1233 1916 1236
rect 1108 1223 1117 1226
rect 1530 1223 1540 1226
rect 1564 1223 1589 1226
rect 1764 1223 1773 1226
rect 1058 1213 1090 1216
rect 1106 1213 1125 1216
rect 1186 1213 1212 1216
rect 1244 1213 1285 1216
rect 1322 1213 1332 1216
rect 1420 1213 1429 1216
rect 1492 1213 1525 1216
rect 1570 1213 1636 1216
rect 1106 1206 1109 1213
rect 122 1203 132 1206
rect 370 1203 381 1206
rect 386 1203 404 1206
rect 476 1203 485 1206
rect 540 1203 557 1206
rect 610 1203 628 1206
rect 642 1203 661 1206
rect 764 1203 789 1206
rect 828 1203 853 1206
rect 908 1203 917 1206
rect 938 1203 965 1206
rect 978 1203 987 1206
rect 1050 1203 1083 1206
rect 1114 1203 1132 1206
rect 1194 1203 1220 1206
rect 1236 1203 1245 1206
rect 1290 1203 1324 1206
rect 1348 1203 1381 1206
rect 1426 1203 1476 1206
rect 1570 1203 1573 1213
rect 1660 1203 1685 1206
rect 378 1196 381 1203
rect 1378 1196 1381 1203
rect 378 1193 389 1196
rect 922 1193 965 1196
rect 1146 1193 1197 1196
rect 1378 1193 1404 1196
rect 1770 1193 1773 1223
rect 1778 1216 1781 1233
rect 1778 1213 1789 1216
rect 1826 1215 1829 1233
rect 1844 1223 1853 1226
rect 1890 1223 1900 1226
rect 2164 1223 2173 1226
rect 2202 1216 2205 1236
rect 2300 1223 2333 1226
rect 2578 1223 2597 1226
rect 2636 1223 2677 1226
rect 3012 1223 3029 1226
rect 3060 1223 3085 1226
rect 2578 1216 2581 1223
rect 1938 1213 1964 1216
rect 2026 1213 2085 1216
rect 2092 1213 2125 1216
rect 2202 1213 2212 1216
rect 2242 1213 2284 1216
rect 2298 1213 2348 1216
rect 2410 1213 2420 1216
rect 2434 1213 2468 1216
rect 2492 1213 2501 1216
rect 2506 1213 2517 1216
rect 2532 1213 2557 1216
rect 2572 1213 2581 1216
rect 2586 1213 2621 1216
rect 2716 1213 2733 1216
rect 2770 1213 2812 1216
rect 2850 1213 2900 1216
rect 2026 1206 2029 1213
rect 1962 1203 1972 1206
rect 1988 1203 2029 1206
rect 2042 1203 2052 1206
rect 2082 1205 2085 1213
rect 2122 1206 2125 1213
rect 2122 1203 2140 1206
rect 2164 1203 2205 1206
rect 2210 1203 2220 1206
rect 2330 1203 2340 1206
rect 2442 1203 2476 1206
rect 2506 1196 2509 1213
rect 2524 1203 2533 1206
rect 2538 1203 2557 1206
rect 2578 1203 2604 1206
rect 2618 1205 2621 1213
rect 2938 1206 2941 1216
rect 2954 1213 2996 1216
rect 3026 1213 3044 1216
rect 2658 1203 2692 1206
rect 2708 1203 2717 1206
rect 2722 1203 2748 1206
rect 2772 1203 2781 1206
rect 2810 1203 2820 1206
rect 2836 1203 2861 1206
rect 2866 1203 2892 1206
rect 2932 1203 2941 1206
rect 2954 1203 2988 1206
rect 3058 1205 3061 1216
rect 3090 1213 3108 1216
rect 3226 1206 3229 1256
rect 3292 1213 3301 1216
rect 3306 1213 3340 1216
rect 3370 1206 3373 1213
rect 3132 1203 3141 1206
rect 3146 1203 3188 1206
rect 3226 1203 3268 1206
rect 3314 1203 3348 1206
rect 3370 1203 3381 1206
rect 2236 1193 2253 1196
rect 2492 1193 2509 1196
rect 2858 1196 2861 1203
rect 2858 1193 2869 1196
rect 1018 1183 1061 1186
rect 3378 1183 3381 1203
rect 38 1167 3434 1173
rect 3290 1153 3317 1156
rect 194 1143 204 1146
rect 370 1143 389 1146
rect 370 1136 373 1143
rect 754 1136 757 1146
rect 2378 1143 2389 1146
rect 2658 1143 2676 1146
rect 90 1133 108 1136
rect 122 1133 156 1136
rect 202 1133 212 1136
rect 274 1133 292 1136
rect 356 1133 373 1136
rect 378 1133 411 1136
rect 428 1133 461 1136
rect 546 1133 563 1136
rect 580 1133 629 1136
rect 660 1133 701 1136
rect 732 1133 741 1136
rect 754 1133 771 1136
rect 458 1126 461 1133
rect 124 1123 141 1126
rect 234 1123 269 1126
rect 300 1123 309 1126
rect 364 1123 389 1126
rect 458 1123 476 1126
rect 524 1123 541 1126
rect 588 1123 635 1126
rect 668 1123 685 1126
rect 690 1123 708 1126
rect 746 1123 778 1126
rect 782 1123 797 1126
rect 802 1116 805 1136
rect 810 1133 820 1136
rect 810 1123 828 1126
rect 308 1113 325 1116
rect 794 1113 805 1116
rect 834 1115 837 1136
rect 842 1133 852 1136
rect 882 1133 892 1136
rect 970 1133 980 1136
rect 1050 1133 1092 1136
rect 1130 1133 1164 1136
rect 1194 1133 1236 1136
rect 1274 1133 1308 1136
rect 1322 1133 1380 1136
rect 1404 1133 1429 1136
rect 1476 1133 1493 1136
rect 1540 1133 1589 1136
rect 1620 1133 1629 1136
rect 1634 1133 1692 1136
rect 1722 1133 1764 1136
rect 1810 1133 1836 1136
rect 1922 1133 1940 1136
rect 2034 1133 2068 1136
rect 2130 1133 2140 1136
rect 2226 1133 2260 1136
rect 866 1123 900 1126
rect 930 1123 948 1126
rect 962 1123 988 1126
rect 1018 1123 1061 1126
rect 1162 1123 1172 1126
rect 1218 1123 1228 1126
rect 1260 1123 1316 1126
rect 1442 1123 1460 1126
rect 1570 1123 1596 1126
rect 1634 1123 1709 1126
rect 1722 1123 1756 1126
rect 1780 1123 1797 1126
rect 1844 1123 1869 1126
rect 908 1113 925 1116
rect 996 1113 1005 1116
rect 1002 1093 1005 1113
rect 1018 1103 1021 1123
rect 1922 1116 1925 1133
rect 2306 1126 2309 1136
rect 2354 1133 2364 1136
rect 2386 1126 2389 1143
rect 2866 1136 2869 1146
rect 3076 1143 3117 1146
rect 3170 1136 3173 1146
rect 2452 1133 2517 1136
rect 2562 1133 2580 1136
rect 2658 1133 2684 1136
rect 2690 1133 2708 1136
rect 2850 1133 2892 1136
rect 2914 1133 2925 1136
rect 2930 1133 2948 1136
rect 2986 1133 2996 1136
rect 3082 1133 3140 1136
rect 3156 1133 3173 1136
rect 3354 1133 3364 1136
rect 2922 1126 2925 1133
rect 1938 1123 1948 1126
rect 2026 1123 2060 1126
rect 2098 1123 2148 1126
rect 2196 1123 2237 1126
rect 2242 1123 2252 1126
rect 2284 1123 2309 1126
rect 2372 1123 2381 1126
rect 2386 1123 2428 1126
rect 2506 1123 2516 1126
rect 2548 1123 2557 1126
rect 2610 1123 2644 1126
rect 2698 1123 2788 1126
rect 2922 1123 2956 1126
rect 3034 1123 3052 1126
rect 3076 1123 3085 1126
rect 3178 1123 3228 1126
rect 3260 1123 3301 1126
rect 3322 1123 3332 1126
rect 3338 1123 3348 1126
rect 3354 1123 3372 1126
rect 2234 1116 2237 1123
rect 1036 1113 1045 1116
rect 1180 1113 1221 1116
rect 1324 1113 1365 1116
rect 1476 1113 1525 1116
rect 1916 1113 1925 1116
rect 2020 1113 2037 1116
rect 2234 1113 2245 1116
rect 1042 1083 1045 1113
rect 1850 1103 1908 1106
rect 1986 1103 2012 1106
rect 14 1067 3458 1073
rect 730 1053 749 1056
rect 818 1043 837 1046
rect 818 1033 829 1036
rect 834 1026 837 1043
rect 244 1023 293 1026
rect 644 1023 669 1026
rect 818 1023 837 1026
rect 898 1023 901 1046
rect 3066 1043 3077 1046
rect 1794 1033 1845 1036
rect 1188 1023 1197 1026
rect 1644 1023 1653 1026
rect 186 1013 204 1016
rect 218 1013 277 1016
rect 316 1013 325 1016
rect 412 1013 445 1016
rect 450 1006 453 1015
rect 498 1013 524 1016
rect 594 1013 628 1016
rect 642 1013 692 1016
rect 718 1013 773 1016
rect 812 1013 845 1016
rect 946 1013 956 1016
rect 988 1013 1013 1016
rect 1018 1013 1036 1016
rect 1068 1013 1101 1016
rect 1138 1013 1172 1016
rect 1194 1013 1244 1016
rect 1250 1013 1284 1016
rect 1396 1013 1429 1016
rect 1516 1013 1533 1016
rect 1602 1013 1636 1016
rect 1642 1013 1676 1016
rect 1746 1013 1788 1016
rect 1842 1015 1845 1033
rect 2978 1033 3013 1036
rect 1924 1023 1949 1026
rect 2236 1023 2285 1026
rect 1866 1013 1908 1016
rect 1972 1013 2012 1016
rect 2068 1013 2085 1016
rect 2124 1013 2133 1016
rect 2146 1013 2212 1016
rect 2258 1013 2292 1016
rect 2316 1013 2333 1016
rect 2338 1013 2364 1016
rect 2420 1013 2453 1016
rect 498 1006 501 1013
rect 210 1003 228 1006
rect 418 1003 453 1006
rect 476 1003 501 1006
rect 530 1003 563 1006
rect 588 1003 613 1006
rect 650 1003 684 1006
rect 698 1003 708 1006
rect 778 1003 788 1006
rect 804 1003 845 1006
rect 980 1003 1005 1006
rect 1194 1003 1197 1013
rect 1308 1003 1325 1006
rect 1338 1003 1388 1006
rect 1410 1003 1436 1006
rect 1450 1003 1508 1006
rect 1546 1003 1556 1006
rect 1682 1003 1732 1006
rect 1930 1003 1964 1006
rect 2034 1003 2060 1006
rect 2074 1003 2100 1006
rect 2154 1003 2204 1006
rect 2234 1003 2300 1006
rect 2338 1003 2356 1006
rect 2386 1003 2412 1006
rect 2418 1003 2460 1006
rect 2530 1003 2564 1006
rect 2338 996 2341 1003
rect 2570 996 2573 1015
rect 2604 1013 2661 1016
rect 2684 1013 2708 1016
rect 2828 1013 2837 1016
rect 2876 1013 2901 1016
rect 2922 1013 2932 1016
rect 2964 1013 2973 1016
rect 2834 1006 2837 1013
rect 2978 1006 2981 1033
rect 3044 1023 3069 1026
rect 3074 1016 3077 1043
rect 3106 1016 3109 1036
rect 3172 1023 3205 1026
rect 3228 1023 3261 1026
rect 3348 1023 3397 1026
rect 3002 1013 3028 1016
rect 3066 1013 3093 1016
rect 3100 1013 3109 1016
rect 3220 1013 3229 1016
rect 3258 1013 3261 1023
rect 3298 1013 3340 1016
rect 2586 1003 2596 1006
rect 2626 1003 2676 1006
rect 2682 1003 2700 1006
rect 2730 1003 2748 1006
rect 2778 1003 2820 1006
rect 2834 1003 2860 1006
rect 2914 1003 2940 1006
rect 2970 1003 2981 1006
rect 2994 1003 3020 1006
rect 3044 1003 3085 1006
rect 3090 1005 3093 1013
rect 3242 1003 3276 1006
rect 3314 1003 3332 1006
rect 3394 1003 3397 1023
rect 2586 996 2589 1003
rect 834 993 852 996
rect 1322 993 1380 996
rect 1482 993 1500 996
rect 2316 993 2341 996
rect 2418 993 2452 996
rect 2546 993 2556 996
rect 2570 993 2589 996
rect 2650 993 2668 996
rect 2770 993 2812 996
rect 3066 993 3085 996
rect 818 983 837 986
rect 906 983 933 986
rect 38 967 3434 973
rect 618 953 637 956
rect 346 936 349 946
rect 906 943 916 946
rect 1050 943 1061 946
rect 130 933 140 936
rect 194 933 204 936
rect 346 933 388 936
rect 402 926 405 936
rect 546 933 588 936
rect 714 933 740 936
rect 770 933 811 936
rect 818 933 836 936
rect 850 926 853 936
rect 858 933 884 936
rect 924 933 957 936
rect 970 933 980 936
rect 954 926 957 933
rect 1002 926 1005 934
rect 1018 933 1036 936
rect 1050 926 1053 943
rect 1122 936 1125 956
rect 1130 953 1149 956
rect 1058 933 1090 936
rect 1108 933 1125 936
rect 1146 936 1149 953
rect 1146 933 1164 936
rect 1244 933 1277 936
rect 1298 926 1301 946
rect 1378 943 1428 946
rect 1522 943 1540 946
rect 2306 943 2324 946
rect 2498 943 2509 946
rect 1364 933 1373 936
rect 1426 933 1436 936
rect 1450 933 1484 936
rect 1490 933 1548 936
rect 1554 933 1596 936
rect 1626 933 1660 936
rect 1682 933 1716 936
rect 2026 933 2052 936
rect 2122 933 2132 936
rect 2156 933 2165 936
rect 2236 933 2269 936
rect 2332 933 2357 936
rect 2418 933 2429 936
rect 2434 933 2453 936
rect 148 923 165 926
rect 330 923 340 926
rect 346 923 405 926
rect 100 913 109 916
rect 124 913 133 916
rect 156 913 189 916
rect 228 913 237 916
rect 266 913 309 916
rect 452 913 461 916
rect 506 906 509 925
rect 540 923 573 926
rect 98 903 116 906
rect 226 903 244 906
rect 258 903 316 906
rect 490 903 509 906
rect 546 903 549 923
rect 626 913 644 916
rect 650 906 653 925
rect 690 923 708 926
rect 850 923 892 926
rect 954 923 987 926
rect 1002 923 1021 926
rect 1044 923 1053 926
rect 1074 923 1083 926
rect 1194 923 1220 926
rect 1252 923 1261 926
rect 1274 923 1324 926
rect 1492 923 1533 926
rect 1578 923 1604 926
rect 1668 923 1685 926
rect 1698 923 1724 926
rect 1746 923 1804 926
rect 1818 923 1844 926
rect 1908 923 1941 926
rect 2034 923 2060 926
rect 2154 923 2212 926
rect 2250 923 2292 926
rect 2354 923 2357 933
rect 2378 923 2388 926
rect 716 913 725 916
rect 1004 913 1013 916
rect 634 903 653 906
rect 682 903 701 906
rect 722 903 725 913
rect 1018 903 1021 923
rect 1074 916 1077 923
rect 1050 913 1077 916
rect 1122 903 1157 906
rect 850 893 869 896
rect 946 893 973 896
rect 1258 893 1261 923
rect 1578 913 1581 923
rect 1612 913 1637 916
rect 1676 913 1709 916
rect 1732 913 1741 916
rect 1820 913 1829 916
rect 1964 913 1989 916
rect 2300 913 2309 916
rect 2098 903 2125 906
rect 2426 896 2429 933
rect 2434 923 2476 926
rect 2498 916 2501 943
rect 2682 936 2685 946
rect 2762 943 2804 946
rect 2556 933 2597 936
rect 2682 933 2716 936
rect 2762 933 2812 936
rect 2986 933 3004 936
rect 3034 933 3044 936
rect 3068 933 3117 936
rect 2506 923 2532 926
rect 2562 923 2581 926
rect 2642 923 2652 926
rect 2740 923 2749 926
rect 2764 923 2805 926
rect 2498 913 2509 916
rect 2834 913 2844 916
rect 2882 913 2908 916
rect 2914 906 2917 925
rect 2954 923 2964 926
rect 3082 923 3124 926
rect 3146 923 3149 934
rect 3226 933 3252 936
rect 3156 923 3189 926
rect 3218 923 3244 926
rect 3276 923 3285 926
rect 3290 923 3340 926
rect 3354 923 3364 926
rect 3186 913 3189 923
rect 3282 916 3285 923
rect 3282 913 3301 916
rect 2826 903 2860 906
rect 2874 903 2917 906
rect 1690 893 1709 896
rect 2426 893 2437 896
rect 14 867 3458 873
rect 1210 853 1237 856
rect 114 833 133 836
rect 338 826 341 846
rect 108 823 141 826
rect 156 823 189 826
rect 330 823 341 826
rect 516 823 557 826
rect 596 823 605 826
rect 820 823 845 826
rect 1092 823 1133 826
rect 1148 823 1157 826
rect 1204 823 1221 826
rect 602 816 605 823
rect 1386 816 1389 826
rect 1666 823 1677 826
rect 1820 823 1853 826
rect 66 813 100 816
rect 148 813 173 816
rect 234 813 277 816
rect 316 813 325 816
rect 412 813 437 816
rect 468 813 485 816
rect 602 813 613 816
rect 274 806 277 813
rect 66 803 92 806
rect 130 803 140 806
rect 178 803 204 806
rect 220 803 269 806
rect 274 803 292 806
rect 434 803 452 806
rect 620 803 653 806
rect 658 783 661 816
rect 700 813 709 816
rect 818 813 837 816
rect 906 813 916 816
rect 970 813 1004 816
rect 1066 813 1076 816
rect 1114 813 1125 816
rect 1140 813 1149 816
rect 1250 813 1268 816
rect 1356 813 1365 816
rect 1386 813 1396 816
rect 1428 813 1477 816
rect 706 805 709 813
rect 740 803 796 806
rect 834 783 837 813
rect 1122 806 1125 813
rect 1474 806 1477 813
rect 1506 813 1532 816
rect 1506 806 1509 813
rect 898 803 924 806
rect 962 803 996 806
rect 1020 803 1061 806
rect 1092 803 1117 806
rect 1122 803 1132 806
rect 1204 803 1237 806
rect 1292 803 1301 806
rect 1348 803 1389 806
rect 1420 803 1469 806
rect 1474 803 1492 806
rect 1498 803 1509 806
rect 1562 806 1565 815
rect 1570 813 1620 816
rect 1652 813 1669 816
rect 1674 806 1677 823
rect 1700 813 1741 816
rect 1756 813 1797 816
rect 1850 806 1853 823
rect 2034 816 2037 825
rect 1972 813 1997 816
rect 2034 813 2045 816
rect 2052 813 2108 816
rect 2178 813 2212 816
rect 2218 813 2228 816
rect 2282 813 2316 816
rect 2436 813 2445 816
rect 2466 806 2469 836
rect 2850 833 2876 836
rect 3002 833 3020 836
rect 2500 823 2533 826
rect 2890 823 2916 826
rect 2940 823 2949 826
rect 3028 823 3053 826
rect 3084 823 3117 826
rect 3380 823 3405 826
rect 3050 816 3053 823
rect 2482 813 2492 816
rect 2514 813 2525 816
rect 2556 813 2581 816
rect 2522 806 2525 813
rect 2690 806 2693 815
rect 2722 813 2756 816
rect 2946 813 2988 816
rect 3050 813 3068 816
rect 3098 813 3132 816
rect 3194 813 3204 816
rect 3258 813 3268 816
rect 3314 813 3348 816
rect 3362 813 3372 816
rect 1562 803 1581 806
rect 1602 803 1628 806
rect 1674 803 1692 806
rect 1722 803 1748 806
rect 1770 803 1796 806
rect 1850 803 1861 806
rect 1884 803 1933 806
rect 1964 803 1989 806
rect 2124 803 2133 806
rect 2140 803 2149 806
rect 2154 803 2204 806
rect 2234 803 2252 806
rect 2378 803 2428 806
rect 2434 803 2444 806
rect 2466 803 2484 806
rect 2522 803 2548 806
rect 2594 803 2604 806
rect 2668 803 2693 806
rect 3050 803 3060 806
rect 3106 803 3124 806
rect 3156 803 3189 806
rect 3228 803 3253 806
rect 3266 803 3276 806
rect 3322 803 3340 806
rect 2146 796 2149 803
rect 1722 793 1740 796
rect 2146 793 2173 796
rect 2394 793 2420 796
rect 2506 793 2540 796
rect 2554 793 2580 796
rect 2634 793 2660 796
rect 2716 793 2725 796
rect 38 767 3434 773
rect 90 733 100 736
rect 170 726 173 756
rect 602 736 605 745
rect 1330 743 1364 746
rect 1482 743 1524 746
rect 1546 743 1564 746
rect 1786 743 1796 746
rect 1898 743 1948 746
rect 2114 743 2133 746
rect 2370 743 2380 746
rect 2394 743 2436 746
rect 2810 743 2836 746
rect 3178 743 3188 746
rect 202 733 213 736
rect 218 733 236 736
rect 252 733 285 736
rect 354 733 364 736
rect 386 733 404 736
rect 442 733 484 736
rect 506 733 516 736
rect 596 733 605 736
rect 650 733 668 736
rect 788 733 820 736
rect 844 733 853 736
rect 858 733 892 736
rect 908 733 956 736
rect 1002 733 1012 736
rect 1042 733 1068 736
rect 1098 733 1117 736
rect 1138 733 1148 736
rect 1250 734 1260 736
rect 1250 733 1261 734
rect 1274 733 1324 736
rect 1338 733 1372 736
rect 1402 733 1444 736
rect 1460 733 1501 736
rect 1514 733 1532 736
rect 1554 733 1572 736
rect 1730 733 1756 736
rect 1810 733 1868 736
rect 1884 733 1893 736
rect 1938 733 2020 736
rect 2036 733 2101 736
rect 2108 733 2117 736
rect 66 723 92 726
rect 124 723 133 726
rect 66 713 69 723
rect 130 696 133 723
rect 164 713 173 716
rect 202 706 205 733
rect 210 723 228 726
rect 306 706 309 725
rect 354 723 372 726
rect 378 723 396 726
rect 466 723 476 726
rect 506 725 509 733
rect 1258 726 1261 733
rect 2154 726 2157 734
rect 2180 733 2189 736
rect 2194 733 2220 736
rect 2276 733 2293 736
rect 2354 733 2388 736
rect 2402 733 2444 736
rect 2458 733 2469 736
rect 2650 733 2660 736
rect 2690 733 2740 736
rect 2788 733 2805 736
rect 2850 733 2869 736
rect 2930 733 2940 736
rect 2458 726 2461 733
rect 514 723 524 726
rect 562 723 580 726
rect 708 723 757 726
rect 818 723 828 726
rect 874 723 884 726
rect 988 723 997 726
rect 1002 723 1020 726
rect 1098 723 1132 726
rect 1156 723 1165 726
rect 1220 723 1261 726
rect 1268 723 1317 726
rect 1332 723 1365 726
rect 1540 723 1565 726
rect 1716 723 1725 726
rect 1764 723 1773 726
rect 1812 723 1853 726
rect 1892 723 1941 726
rect 1978 723 2012 726
rect 2044 723 2061 726
rect 2116 723 2157 726
rect 2284 723 2309 726
rect 2340 723 2365 726
rect 2452 723 2461 726
rect 2466 723 2500 726
rect 2530 723 2580 726
rect 2618 723 2644 726
rect 2650 723 2668 726
rect 2748 723 2772 726
rect 2866 716 2869 733
rect 3042 726 3045 734
rect 3106 733 3172 736
rect 3218 733 3292 736
rect 380 713 389 716
rect 844 713 861 716
rect 1028 713 1053 716
rect 1644 713 1653 716
rect 2348 713 2373 716
rect 2516 713 2565 716
rect 2684 713 2709 716
rect 2788 713 2829 716
rect 138 703 165 706
rect 202 703 221 706
rect 290 703 309 706
rect 130 693 141 696
rect 386 683 389 713
rect 2858 706 2861 716
rect 2866 713 2876 716
rect 2882 706 2885 725
rect 2906 723 2948 726
rect 3034 723 3045 726
rect 3180 723 3189 726
rect 3226 723 3284 726
rect 3034 716 3037 723
rect 2900 713 2909 716
rect 2954 713 2980 716
rect 3004 713 3037 716
rect 3100 713 3157 716
rect 1586 703 1660 706
rect 2858 703 2885 706
rect 2978 703 2996 706
rect 14 667 3458 673
rect 426 633 461 636
rect 506 633 532 636
rect 634 633 661 636
rect 108 623 117 626
rect 266 623 277 626
rect 332 623 349 626
rect 266 616 269 623
rect 426 616 429 633
rect 434 623 452 626
rect 476 623 485 626
rect 498 623 516 626
rect 172 613 213 616
rect 252 613 269 616
rect 274 613 300 616
rect 306 613 324 616
rect 330 613 388 616
rect 420 613 429 616
rect 594 613 628 616
rect 658 615 661 633
rect 874 626 877 636
rect 1578 633 1612 636
rect 1874 626 1877 636
rect 2378 633 2404 636
rect 2594 633 2620 636
rect 844 623 877 626
rect 892 623 925 626
rect 1052 623 1069 626
rect 1220 623 1237 626
rect 1444 623 1453 626
rect 1620 623 1637 626
rect 1740 623 1789 626
rect 1868 623 1877 626
rect 2100 623 2133 626
rect 780 613 813 616
rect 858 613 884 616
rect 890 613 948 616
rect 1002 613 1036 616
rect 1108 613 1117 616
rect 1164 613 1189 616
rect 1194 613 1204 616
rect 1226 613 1277 616
rect 1346 613 1356 616
rect 1394 613 1428 616
rect 1442 613 1500 616
rect 1626 613 1668 616
rect 1738 613 1773 616
rect 1812 613 1837 616
rect 1842 613 1852 616
rect 1866 613 1924 616
rect 1956 613 2013 616
rect 2226 613 2268 616
rect 2292 613 2309 616
rect 210 606 213 613
rect 274 606 277 613
rect 130 603 148 606
rect 164 603 197 606
rect 210 603 221 606
rect 244 603 277 606
rect 378 603 396 606
rect 724 603 733 606
rect 772 603 781 606
rect 810 603 820 606
rect 930 603 940 606
rect 978 603 1028 606
rect 1052 603 1061 606
rect 1066 603 1083 606
rect 1114 603 1140 606
rect 1220 603 1269 606
rect 1274 605 1277 613
rect 1308 603 1317 606
rect 1322 603 1348 606
rect 1378 603 1420 606
rect 1490 603 1508 606
rect 1626 603 1660 606
rect 1682 603 1716 606
rect 1738 605 1741 613
rect 2378 606 2381 633
rect 2412 623 2437 626
rect 2484 623 2501 626
rect 3188 623 3221 626
rect 3252 623 3269 626
rect 3314 623 3333 626
rect 2442 613 2468 616
rect 2514 613 2532 616
rect 2634 613 2676 616
rect 2826 613 2852 616
rect 3052 613 3061 616
rect 3068 613 3101 616
rect 3132 613 3141 616
rect 3162 613 3237 616
rect 3244 613 3269 616
rect 3356 613 3365 616
rect 3380 613 3397 616
rect 1746 603 1804 606
rect 1810 603 1844 606
rect 1868 603 1877 606
rect 1890 603 1932 606
rect 2036 603 2061 606
rect 2106 603 2148 606
rect 2170 603 2204 606
rect 2226 603 2260 606
rect 2284 603 2301 606
rect 2364 603 2381 606
rect 2418 603 2460 606
rect 2484 603 2493 606
rect 2522 603 2540 606
rect 2642 603 2684 606
rect 2700 603 2741 606
rect 2754 603 2773 606
rect 2914 603 2948 606
rect 2954 603 2997 606
rect 3186 603 3236 606
rect 3250 603 3284 606
rect 682 593 716 596
rect 2220 593 2253 596
rect 2714 593 2740 596
rect 2914 593 2940 596
rect 3074 593 3116 596
rect 38 567 3434 573
rect 730 536 733 545
rect 1274 543 1324 546
rect 1370 543 1396 546
rect 1650 543 1677 546
rect 2170 543 2205 546
rect 1650 536 1653 543
rect 162 533 204 536
rect 220 533 285 536
rect 322 533 388 536
rect 650 533 700 536
rect 724 533 733 536
rect 810 533 820 536
rect 858 533 876 536
rect 930 533 940 536
rect 1170 533 1188 536
rect 1298 533 1332 536
rect 1404 533 1413 536
rect 1602 533 1612 536
rect 1636 533 1653 536
rect 1658 533 1708 536
rect 1724 533 1733 536
rect 1738 533 1788 536
rect 2042 533 2060 536
rect 2148 533 2165 536
rect 2178 533 2212 536
rect 2226 533 2269 536
rect 2338 533 2348 536
rect 66 523 100 526
rect 122 523 140 526
rect 178 523 196 526
rect 228 523 253 526
rect 258 523 292 526
rect 324 523 341 526
rect 386 523 396 526
rect 420 523 469 526
rect 532 523 589 526
rect 626 523 701 526
rect 756 523 773 526
rect 858 523 884 526
rect 948 523 965 526
rect 148 513 189 516
rect 562 513 596 516
rect 954 513 972 516
rect 1018 513 1052 516
rect 1082 513 1124 516
rect 1130 506 1133 525
rect 1170 516 1173 533
rect 1412 523 1445 526
rect 1594 523 1620 526
rect 1746 523 1796 526
rect 1818 523 1852 526
rect 1866 523 1908 526
rect 1940 523 1957 526
rect 2026 523 2068 526
rect 2098 523 2124 526
rect 2156 523 2205 526
rect 2220 523 2261 526
rect 2266 525 2269 533
rect 2370 526 2373 556
rect 2420 533 2437 536
rect 2458 533 2484 536
rect 2650 533 2676 536
rect 2778 533 2828 536
rect 2850 526 2853 535
rect 2938 526 2941 536
rect 3042 526 3045 545
rect 3058 543 3076 546
rect 3052 533 3069 536
rect 3122 533 3140 536
rect 3122 526 3125 533
rect 2356 523 2373 526
rect 2378 523 2396 526
rect 2428 523 2461 526
rect 2492 523 2501 526
rect 2578 523 2612 526
rect 2634 523 2644 526
rect 2690 523 2732 526
rect 2754 523 2764 526
rect 2850 523 2861 526
rect 2868 523 2877 526
rect 2932 523 2941 526
rect 2946 523 2964 526
rect 2988 523 3045 526
rect 3092 523 3125 526
rect 3170 523 3196 526
rect 3242 523 3284 526
rect 3316 523 3349 526
rect 1594 516 1597 523
rect 1148 513 1173 516
rect 1226 513 1236 516
rect 1260 513 1269 516
rect 1484 513 1533 516
rect 1538 506 1541 515
rect 1564 513 1597 516
rect 1636 513 1677 516
rect 1746 513 1749 523
rect 1804 513 1845 516
rect 1860 513 1901 516
rect 2076 513 2117 516
rect 1002 503 1068 506
rect 1114 503 1133 506
rect 1202 503 1252 506
rect 1426 503 1476 506
rect 1506 503 1541 506
rect 3346 506 3349 523
rect 3346 503 3372 506
rect 1002 493 1005 503
rect 14 467 3458 473
rect 362 426 365 436
rect 698 433 724 436
rect 2090 433 2124 436
rect 3338 433 3364 436
rect 324 423 365 426
rect 588 423 621 426
rect 858 416 861 426
rect 1492 423 1509 426
rect 1564 423 1573 426
rect 1692 423 1701 426
rect 1882 423 1917 426
rect 2098 423 2108 426
rect 2132 423 2165 426
rect 2972 423 3021 426
rect 3068 423 3101 426
rect 3276 423 3309 426
rect 3338 423 3348 426
rect 3372 423 3381 426
rect 1882 416 1885 423
rect 124 413 180 416
rect 212 413 245 416
rect 266 413 292 416
rect 298 413 365 416
rect 372 413 381 416
rect 426 413 452 416
rect 508 413 517 416
rect 524 413 572 416
rect 738 413 764 416
rect 836 413 845 416
rect 858 413 868 416
rect 906 413 964 416
rect 1002 413 1012 416
rect 1034 413 1068 416
rect 1140 413 1157 416
rect 1188 413 1237 416
rect 116 403 149 406
rect 204 403 237 406
rect 242 405 245 413
rect 258 403 284 406
rect 770 403 781 406
rect 786 403 820 406
rect 850 403 876 406
rect 930 403 956 406
rect 980 403 997 406
rect 1084 403 1109 406
rect 1234 405 1237 413
rect 1290 413 1332 416
rect 1338 413 1356 416
rect 1466 413 1476 416
rect 1610 413 1620 416
rect 1684 413 1741 416
rect 1828 413 1861 416
rect 1868 413 1885 416
rect 1890 413 1924 416
rect 1946 413 1981 416
rect 2194 413 2213 416
rect 2284 413 2293 416
rect 2322 413 2332 416
rect 2356 413 2397 416
rect 2426 413 2437 416
rect 2530 413 2556 416
rect 2692 413 2716 416
rect 2730 413 2780 416
rect 2818 413 2836 416
rect 2868 413 2893 416
rect 2940 413 2949 416
rect 2994 413 3036 416
rect 3042 413 3052 416
rect 3140 413 3181 416
rect 3234 413 3268 416
rect 3274 413 3324 416
rect 1290 406 1293 413
rect 2210 406 2213 413
rect 1268 403 1293 406
rect 1338 403 1348 406
rect 1378 403 1396 406
rect 1450 403 1468 406
rect 1498 403 1540 406
rect 1564 403 1573 406
rect 1594 403 1612 406
rect 1650 403 1676 406
rect 1764 403 1781 406
rect 1786 403 1860 406
rect 1930 403 1948 406
rect 2196 403 2205 406
rect 2210 403 2260 406
rect 2330 403 2340 406
rect 2426 405 2429 413
rect 2434 403 2484 406
rect 2500 403 2517 406
rect 2538 403 2548 406
rect 2610 403 2620 406
rect 2732 403 2773 406
rect 2860 403 2909 406
rect 2914 403 2948 406
rect 3002 403 3028 406
rect 3132 403 3157 406
rect 3220 403 3253 406
rect 146 383 149 403
rect 778 396 781 403
rect 1106 396 1109 403
rect 458 393 492 396
rect 778 393 812 396
rect 1106 393 1116 396
rect 2434 393 2437 403
rect 2906 393 2924 396
rect 38 367 3434 373
rect 2348 343 2357 346
rect 66 333 100 336
rect 130 333 140 336
rect 162 333 196 336
rect 226 333 236 336
rect 266 333 292 336
rect 490 333 500 336
rect 266 326 269 333
rect 522 326 525 334
rect 530 333 548 336
rect 572 333 621 336
rect 700 333 709 336
rect 770 333 780 336
rect 818 333 828 336
rect 906 333 948 336
rect 978 333 1028 336
rect 1058 333 1077 336
rect 1108 333 1125 336
rect 1410 333 1428 336
rect 1442 333 1468 336
rect 1554 333 1572 336
rect 1596 333 1605 336
rect 1730 333 1748 336
rect 1786 333 1812 336
rect 1828 333 1893 336
rect 1986 333 2004 336
rect 2066 333 2076 336
rect 2100 333 2109 336
rect 2186 333 2204 336
rect 2322 333 2332 336
rect 2434 333 2476 336
rect 2506 333 2548 336
rect 2930 333 2948 336
rect 3082 333 3092 336
rect 3194 333 3212 336
rect 3258 333 3292 336
rect 3308 333 3341 336
rect 1058 326 1061 333
rect 130 323 148 326
rect 186 323 204 326
rect 226 323 244 326
rect 260 323 269 326
rect 322 323 332 326
rect 482 323 508 326
rect 522 323 549 326
rect 610 323 620 326
rect 652 323 669 326
rect 674 323 684 326
rect 698 323 709 326
rect 770 323 788 326
rect 810 323 836 326
rect 914 323 940 326
rect 978 323 1020 326
rect 1052 323 1061 326
rect 1066 323 1092 326
rect 1114 323 1156 326
rect 1364 323 1413 326
rect 1418 323 1436 326
rect 130 313 133 323
rect 156 313 197 316
rect 266 313 269 323
rect 706 316 709 323
rect 1410 316 1413 323
rect 346 313 396 316
rect 452 313 461 316
rect 572 313 597 316
rect 706 313 740 316
rect 852 313 861 316
rect 900 313 909 316
rect 1162 313 1180 316
rect 1204 313 1213 316
rect 1244 313 1253 316
rect 1268 313 1277 316
rect 1410 313 1429 316
rect 1442 315 1445 333
rect 1786 326 1789 333
rect 1756 323 1797 326
rect 1948 323 2005 326
rect 1596 313 1645 316
rect 1924 313 1933 316
rect 2100 313 2149 316
rect 2162 306 2165 325
rect 2186 323 2212 326
rect 2290 323 2324 326
rect 2180 313 2197 316
rect 2234 313 2260 316
rect 2284 313 2301 316
rect 2402 306 2405 325
rect 2426 323 2468 326
rect 2562 323 2572 326
rect 2578 323 2636 326
rect 2650 323 2668 326
rect 2682 323 2708 326
rect 2714 323 2748 326
rect 2938 323 2956 326
rect 2802 313 2836 316
rect 2988 313 3005 316
rect 3018 313 3044 316
rect 3114 313 3156 316
rect 3162 306 3165 325
rect 3202 323 3269 326
rect 3228 313 3253 316
rect 3356 313 3365 316
rect 362 303 412 306
rect 426 303 444 306
rect 1170 303 1196 306
rect 1210 303 1260 306
rect 2106 303 2165 306
rect 2250 303 2276 306
rect 2386 303 2405 306
rect 2786 303 2852 306
rect 2994 303 3060 306
rect 3106 303 3165 306
rect 3322 303 3372 306
rect 14 267 3458 273
rect 162 233 204 236
rect 226 233 268 236
rect 146 223 188 226
rect 252 223 261 226
rect 428 223 445 226
rect 500 223 525 226
rect 794 216 797 236
rect 1106 233 1172 236
rect 1250 233 1260 236
rect 2274 233 2324 236
rect 906 223 925 226
rect 1106 223 1165 226
rect 1180 223 1197 226
rect 1202 223 1244 226
rect 1268 223 1277 226
rect 1466 223 1501 226
rect 1516 223 1533 226
rect 906 216 909 223
rect 1466 216 1469 223
rect 1626 216 1629 226
rect 1780 223 1821 226
rect 1978 223 2005 226
rect 2036 223 2045 226
rect 2066 223 2092 226
rect 2116 223 2149 226
rect 2308 223 2317 226
rect 2332 223 2341 226
rect 2346 223 2372 226
rect 2556 223 2565 226
rect 2660 223 2685 226
rect 132 213 173 216
rect 282 213 340 216
rect 372 213 413 216
rect 420 213 437 216
rect 450 213 484 216
rect 554 213 604 216
rect 642 213 684 216
rect 706 213 724 216
rect 794 213 804 216
rect 810 213 860 216
rect 892 213 909 216
rect 914 213 956 216
rect 1050 213 1100 216
rect 1306 213 1332 216
rect 1370 213 1469 216
rect 1474 213 1508 216
rect 1554 213 1564 216
rect 1578 213 1636 216
rect 1674 213 1748 216
rect 1754 213 1772 216
rect 1818 213 1821 223
rect 2002 216 2005 223
rect 1826 213 1844 216
rect 1908 213 1949 216
rect 1972 213 1997 216
rect 2002 213 2020 216
rect 1370 206 1373 213
rect 1826 206 1829 213
rect 124 203 181 206
rect 370 203 412 206
rect 466 203 476 206
rect 500 203 525 206
rect 540 203 597 206
rect 602 203 612 206
rect 628 203 661 206
rect 740 203 789 206
rect 842 203 868 206
rect 884 203 909 206
rect 938 203 948 206
rect 1362 203 1373 206
rect 1378 203 1428 206
rect 1514 203 1556 206
rect 1586 203 1644 206
rect 1660 203 1733 206
rect 1754 203 1764 206
rect 1802 203 1829 206
rect 1850 203 1900 206
rect 1930 203 1964 206
rect 1986 203 2012 206
rect 2042 203 2045 223
rect 2146 216 2149 223
rect 2146 213 2164 216
rect 2522 213 2540 216
rect 2554 213 2604 216
rect 2634 213 2644 216
rect 2658 213 2685 216
rect 2690 213 2716 216
rect 2786 213 2812 216
rect 2842 213 2860 216
rect 2866 213 2908 216
rect 2924 213 2957 216
rect 3058 213 3092 216
rect 3130 213 3172 216
rect 3210 213 3260 216
rect 3282 213 3300 216
rect 2682 206 2685 213
rect 3378 206 3381 216
rect 2122 203 2172 206
rect 2194 203 2236 206
rect 2260 203 2301 206
rect 2434 203 2452 206
rect 2468 203 2517 206
rect 2562 203 2596 206
rect 2660 203 2677 206
rect 2682 203 2708 206
rect 2732 203 2741 206
rect 2882 203 2900 206
rect 3170 203 3180 206
rect 3196 203 3229 206
rect 3274 203 3308 206
rect 3324 203 3381 206
rect 522 196 525 203
rect 522 193 532 196
rect 2188 193 2221 196
rect 2738 195 2741 203
rect 38 167 3434 173
rect 1194 143 1221 146
rect 1714 143 1732 146
rect 1194 136 1197 143
rect 2370 136 2373 145
rect 2650 143 2660 146
rect 210 133 221 136
rect 292 133 349 136
rect 378 133 444 136
rect 460 133 485 136
rect 490 133 500 136
rect 628 133 677 136
rect 698 133 749 136
rect 772 133 844 136
rect 866 133 924 136
rect 938 133 956 136
rect 970 133 1028 136
rect 1052 133 1069 136
rect 218 126 221 133
rect 82 123 124 126
rect 138 123 180 126
rect 218 123 268 126
rect 300 123 333 126
rect 338 123 348 126
rect 378 125 381 133
rect 482 126 485 133
rect 386 123 436 126
rect 482 123 508 126
rect 530 123 548 126
rect 586 123 604 126
rect 692 123 741 126
rect 746 125 749 133
rect 1074 126 1077 134
rect 1100 133 1149 136
rect 1180 133 1197 136
rect 1202 133 1244 136
rect 1274 133 1332 136
rect 1370 133 1396 136
rect 1418 133 1460 136
rect 1482 126 1485 134
rect 1490 133 1540 136
rect 1562 126 1565 134
rect 1706 133 1740 136
rect 1746 133 1812 136
rect 2052 133 2061 136
rect 2242 133 2260 136
rect 2348 133 2373 136
rect 2466 133 2484 136
rect 868 123 885 126
rect 932 123 949 126
rect 964 123 1029 126
rect 1050 123 1077 126
rect 1194 123 1236 126
rect 1314 123 1324 126
rect 1386 123 1404 126
rect 1482 123 1541 126
rect 1562 123 1573 126
rect 132 113 173 116
rect 556 113 597 116
rect 940 113 957 116
rect 972 113 1021 116
rect 1052 113 1069 116
rect 1100 113 1141 116
rect 1570 106 1573 123
rect 1578 113 1612 116
rect 1618 106 1621 125
rect 1642 123 1700 126
rect 1706 115 1709 133
rect 1748 123 1789 126
rect 1986 123 2028 126
rect 2082 123 2124 126
rect 2154 123 2172 126
rect 2178 123 2236 126
rect 2242 123 2253 126
rect 2268 123 2317 126
rect 2396 123 2405 126
rect 2410 123 2452 126
rect 2492 123 2517 126
rect 2242 115 2245 123
rect 2514 116 2517 123
rect 2650 116 2653 143
rect 2690 133 2724 136
rect 2786 133 2804 136
rect 2818 133 2844 136
rect 2994 133 3060 136
rect 3196 133 3285 136
rect 2738 123 2756 126
rect 2770 123 2812 126
rect 2818 123 2852 126
rect 2970 123 2988 126
rect 3068 123 3084 126
rect 3204 123 3221 126
rect 3324 123 3341 126
rect 2514 113 2524 116
rect 2570 113 2596 116
rect 2620 113 2653 116
rect 2764 113 2797 116
rect 3100 113 3165 116
rect 1570 103 1621 106
rect 2498 103 2540 106
rect 2554 103 2612 106
rect 2 83 93 86
rect 2 6 5 83
rect 14 67 3458 73
rect 38 37 3434 57
rect 14 13 3458 33
rect 2 3 3013 6
<< metal2 >>
rect 14 13 34 3327
rect 38 37 58 3303
rect 170 3176 173 3246
rect 162 3173 173 3176
rect 218 3176 221 3216
rect 218 3173 229 3176
rect 162 3126 165 3173
rect 186 3133 189 3146
rect 202 3133 221 3136
rect 226 3133 229 3173
rect 250 3143 253 3216
rect 218 3126 221 3133
rect 162 3123 173 3126
rect 90 2956 93 3086
rect 170 3083 173 3123
rect 210 3016 213 3126
rect 218 3123 253 3126
rect 74 2953 93 2956
rect 74 2806 77 2953
rect 130 2943 133 3016
rect 90 2813 93 2936
rect 138 2923 141 2996
rect 170 2906 173 2926
rect 162 2903 173 2906
rect 162 2836 165 2903
rect 194 2896 197 2976
rect 202 2966 205 3016
rect 210 3013 229 3016
rect 210 2986 213 2996
rect 218 2993 221 3006
rect 226 2986 229 2996
rect 210 2983 229 2986
rect 210 2973 213 2983
rect 234 2973 237 3116
rect 202 2963 213 2966
rect 202 2916 205 2936
rect 210 2923 213 2963
rect 218 2926 221 2936
rect 242 2933 245 2946
rect 250 2926 253 3123
rect 258 3106 261 3216
rect 274 3193 277 3206
rect 298 3133 301 3206
rect 314 3133 317 3206
rect 338 3203 341 3216
rect 394 3193 397 3216
rect 258 3103 269 3106
rect 298 3103 301 3116
rect 362 3106 365 3126
rect 354 3103 365 3106
rect 266 3036 269 3103
rect 258 3033 269 3036
rect 258 3013 261 3033
rect 258 2983 261 2996
rect 282 2976 285 3006
rect 306 2993 309 3006
rect 314 3003 317 3036
rect 330 3003 333 3046
rect 354 3026 357 3103
rect 354 3023 365 3026
rect 378 3023 381 3056
rect 394 3033 397 3126
rect 402 3103 405 3126
rect 362 3003 365 3023
rect 402 3003 405 3026
rect 410 3013 413 3216
rect 434 3203 437 3226
rect 466 3183 469 3206
rect 442 3136 445 3146
rect 426 3133 445 3136
rect 466 3126 469 3146
rect 362 2983 365 2996
rect 282 2973 301 2976
rect 218 2923 253 2926
rect 202 2913 221 2916
rect 178 2893 197 2896
rect 162 2833 173 2836
rect 74 2803 93 2806
rect 90 2733 93 2803
rect 114 2746 117 2816
rect 122 2793 125 2806
rect 114 2743 121 2746
rect 118 2696 121 2743
rect 114 2693 121 2696
rect 90 2533 93 2606
rect 114 2383 117 2693
rect 130 2636 133 2816
rect 154 2766 157 2816
rect 170 2813 173 2833
rect 154 2763 165 2766
rect 138 2723 141 2746
rect 162 2686 165 2763
rect 178 2716 181 2893
rect 218 2866 221 2913
rect 234 2906 237 2923
rect 258 2913 261 2936
rect 274 2933 277 2946
rect 298 2923 301 2973
rect 378 2933 381 2946
rect 234 2903 245 2906
rect 218 2863 229 2866
rect 186 2803 189 2826
rect 202 2803 205 2816
rect 226 2813 229 2863
rect 242 2816 245 2903
rect 362 2873 365 2926
rect 402 2923 405 2996
rect 426 2943 429 3116
rect 442 3083 445 3116
rect 450 3053 453 3126
rect 462 3123 469 3126
rect 474 3123 477 3136
rect 450 3013 453 3026
rect 442 2966 445 2986
rect 442 2963 449 2966
rect 446 2886 449 2963
rect 462 2946 465 3123
rect 474 3013 477 3116
rect 490 3043 493 3136
rect 498 3116 501 3256
rect 1786 3246 1789 3276
rect 2386 3253 2413 3256
rect 698 3233 733 3236
rect 514 3133 517 3216
rect 546 3213 549 3226
rect 578 3183 581 3206
rect 602 3146 605 3226
rect 626 3203 629 3216
rect 698 3213 701 3233
rect 714 3223 725 3226
rect 706 3213 725 3216
rect 522 3133 525 3146
rect 602 3143 613 3146
rect 498 3113 509 3116
rect 506 3036 509 3113
rect 562 3106 565 3116
rect 578 3113 581 3136
rect 562 3103 573 3106
rect 570 3036 573 3103
rect 610 3096 613 3143
rect 626 3123 629 3146
rect 666 3106 669 3126
rect 602 3093 613 3096
rect 658 3103 669 3106
rect 498 3033 509 3036
rect 498 2976 501 3033
rect 554 3023 557 3036
rect 570 3033 581 3036
rect 474 2973 501 2976
rect 462 2943 469 2946
rect 442 2883 449 2886
rect 234 2813 245 2816
rect 322 2823 365 2826
rect 322 2813 325 2823
rect 234 2796 237 2813
rect 202 2726 205 2796
rect 218 2793 237 2796
rect 290 2793 293 2806
rect 218 2733 221 2793
rect 202 2723 213 2726
rect 178 2713 197 2716
rect 154 2683 165 2686
rect 154 2656 157 2683
rect 154 2653 165 2656
rect 122 2633 133 2636
rect 122 2476 125 2633
rect 130 2613 133 2626
rect 130 2523 133 2596
rect 162 2566 165 2653
rect 194 2646 197 2713
rect 194 2643 205 2646
rect 178 2603 181 2626
rect 194 2573 197 2616
rect 202 2593 205 2643
rect 154 2563 165 2566
rect 154 2543 157 2563
rect 122 2473 141 2476
rect 138 2376 141 2473
rect 114 2373 141 2376
rect 66 1743 69 1996
rect 66 813 69 1736
rect 74 1593 77 2236
rect 90 2203 93 2336
rect 114 2196 117 2373
rect 170 2366 173 2386
rect 162 2363 173 2366
rect 122 2306 125 2326
rect 162 2316 165 2363
rect 178 2323 181 2536
rect 194 2516 197 2526
rect 210 2523 213 2723
rect 218 2706 221 2726
rect 218 2703 225 2706
rect 222 2636 225 2703
rect 234 2683 237 2793
rect 330 2783 333 2816
rect 346 2813 357 2816
rect 362 2813 365 2823
rect 242 2733 245 2746
rect 242 2663 245 2716
rect 250 2713 253 2736
rect 218 2633 225 2636
rect 218 2613 221 2633
rect 218 2593 221 2606
rect 226 2593 229 2606
rect 250 2546 253 2656
rect 258 2613 261 2726
rect 274 2603 277 2756
rect 306 2733 309 2756
rect 346 2656 349 2813
rect 354 2723 357 2736
rect 306 2653 349 2656
rect 306 2606 309 2653
rect 322 2613 325 2626
rect 306 2603 317 2606
rect 314 2586 317 2603
rect 306 2583 317 2586
rect 242 2543 269 2546
rect 242 2533 245 2543
rect 218 2523 229 2526
rect 234 2516 237 2526
rect 194 2513 237 2516
rect 242 2453 245 2526
rect 250 2493 253 2536
rect 266 2533 269 2543
rect 258 2476 261 2526
rect 254 2473 261 2476
rect 254 2386 257 2473
rect 234 2383 257 2386
rect 234 2336 237 2383
rect 194 2323 197 2336
rect 226 2333 237 2336
rect 162 2313 173 2316
rect 122 2303 133 2306
rect 130 2236 133 2303
rect 122 2233 133 2236
rect 122 2203 125 2233
rect 106 2193 117 2196
rect 82 2133 93 2136
rect 98 2133 101 2156
rect 90 2126 93 2133
rect 106 2126 109 2193
rect 130 2133 133 2216
rect 170 2213 173 2313
rect 226 2276 229 2333
rect 242 2286 245 2326
rect 242 2283 253 2286
rect 226 2273 237 2276
rect 202 2223 229 2226
rect 186 2153 189 2206
rect 90 2123 109 2126
rect 114 2123 125 2126
rect 98 2113 101 2123
rect 114 2096 117 2123
rect 106 2093 117 2096
rect 106 2026 109 2093
rect 106 2023 117 2026
rect 82 1983 85 2006
rect 82 1873 85 1936
rect 90 1923 93 2016
rect 106 1943 109 2006
rect 114 2003 117 2023
rect 98 1933 109 1936
rect 114 1933 117 1956
rect 98 1906 101 1933
rect 94 1903 101 1906
rect 94 1826 97 1903
rect 90 1823 97 1826
rect 82 1696 85 1816
rect 90 1803 93 1823
rect 106 1816 109 1916
rect 114 1913 117 1926
rect 98 1813 109 1816
rect 114 1813 117 1856
rect 98 1733 101 1813
rect 106 1803 117 1806
rect 106 1733 109 1786
rect 114 1733 117 1746
rect 90 1723 109 1726
rect 82 1693 93 1696
rect 74 1443 77 1586
rect 82 1583 85 1686
rect 82 1426 85 1556
rect 90 1536 93 1693
rect 98 1543 101 1716
rect 106 1663 109 1716
rect 106 1613 109 1636
rect 114 1623 117 1706
rect 122 1683 125 2116
rect 130 2023 133 2106
rect 130 1833 133 1936
rect 122 1623 125 1666
rect 114 1613 125 1616
rect 90 1533 109 1536
rect 74 1423 85 1426
rect 90 1513 109 1516
rect 74 1213 77 1423
rect 82 1376 85 1416
rect 90 1413 93 1513
rect 90 1383 93 1406
rect 82 1373 93 1376
rect 82 1333 85 1366
rect 82 1306 85 1326
rect 90 1323 93 1373
rect 82 1303 89 1306
rect 86 1236 89 1303
rect 82 1233 89 1236
rect 74 1163 77 1206
rect 66 723 69 806
rect 66 703 69 716
rect 74 686 77 1156
rect 82 986 85 1233
rect 90 1203 93 1216
rect 90 1133 93 1196
rect 98 1133 101 1496
rect 90 1003 93 1126
rect 98 1113 101 1126
rect 82 983 89 986
rect 86 756 89 983
rect 70 683 77 686
rect 82 753 89 756
rect 98 753 101 1016
rect 106 926 109 1506
rect 114 1493 117 1606
rect 122 1593 125 1606
rect 114 1413 117 1426
rect 122 1403 125 1586
rect 130 1563 133 1826
rect 138 1573 141 2146
rect 170 2143 197 2146
rect 146 2086 149 2106
rect 154 2096 157 2116
rect 154 2093 165 2096
rect 146 2083 157 2086
rect 154 2023 157 2083
rect 162 2033 165 2093
rect 146 1853 149 2016
rect 146 1726 149 1846
rect 154 1733 157 1976
rect 162 1923 165 2026
rect 170 1933 173 2143
rect 178 2133 197 2136
rect 178 2103 181 2133
rect 186 2103 189 2116
rect 178 1933 181 2036
rect 186 1943 189 2026
rect 194 1936 197 2016
rect 186 1933 197 1936
rect 202 1926 205 2223
rect 234 2216 237 2273
rect 250 2216 253 2283
rect 258 2223 261 2236
rect 210 2196 213 2216
rect 234 2213 245 2216
rect 250 2213 261 2216
rect 218 2203 229 2206
rect 234 2203 245 2206
rect 258 2203 261 2213
rect 266 2196 269 2526
rect 282 2523 285 2576
rect 306 2526 309 2583
rect 354 2576 357 2616
rect 362 2603 365 2686
rect 370 2653 373 2806
rect 330 2573 357 2576
rect 330 2533 333 2573
rect 362 2566 365 2596
rect 346 2563 365 2566
rect 306 2523 317 2526
rect 282 2436 285 2456
rect 282 2433 293 2436
rect 290 2366 293 2433
rect 282 2363 293 2366
rect 314 2366 317 2523
rect 338 2403 341 2546
rect 346 2543 349 2563
rect 370 2546 373 2616
rect 378 2566 381 2786
rect 386 2586 389 2816
rect 402 2793 405 2806
rect 418 2783 421 2816
rect 426 2803 429 2826
rect 434 2793 437 2806
rect 418 2753 437 2756
rect 394 2713 397 2726
rect 402 2693 405 2726
rect 410 2683 413 2736
rect 418 2733 421 2753
rect 426 2726 429 2746
rect 434 2733 437 2753
rect 426 2723 437 2726
rect 434 2693 437 2716
rect 442 2706 445 2883
rect 458 2866 461 2926
rect 450 2863 461 2866
rect 450 2813 453 2863
rect 458 2733 461 2816
rect 450 2723 461 2726
rect 466 2713 469 2943
rect 474 2803 477 2973
rect 506 2953 509 3016
rect 514 2983 517 3016
rect 530 2966 533 3006
rect 554 3003 557 3016
rect 562 2966 565 3006
rect 522 2956 525 2966
rect 530 2963 565 2966
rect 570 2963 573 3016
rect 522 2953 533 2956
rect 514 2943 525 2946
rect 482 2933 501 2936
rect 506 2933 517 2936
rect 498 2926 501 2933
rect 490 2893 493 2926
rect 498 2923 509 2926
rect 506 2903 509 2916
rect 474 2733 477 2746
rect 442 2703 449 2706
rect 446 2646 449 2703
rect 474 2663 477 2726
rect 446 2643 453 2646
rect 394 2603 397 2626
rect 402 2623 405 2636
rect 386 2583 397 2586
rect 378 2563 385 2566
rect 362 2543 373 2546
rect 362 2526 365 2543
rect 346 2523 365 2526
rect 370 2506 373 2536
rect 366 2503 373 2506
rect 366 2436 369 2503
rect 382 2496 385 2563
rect 378 2493 385 2496
rect 366 2433 373 2436
rect 370 2413 373 2433
rect 378 2376 381 2493
rect 394 2466 397 2583
rect 418 2553 421 2616
rect 450 2596 453 2643
rect 466 2613 469 2626
rect 442 2593 453 2596
rect 442 2546 445 2593
rect 482 2556 485 2856
rect 490 2803 493 2826
rect 498 2813 501 2876
rect 490 2736 493 2786
rect 522 2746 525 2943
rect 530 2853 533 2953
rect 538 2933 541 2963
rect 538 2756 541 2816
rect 554 2813 557 2926
rect 562 2806 565 2836
rect 570 2813 573 2956
rect 578 2933 581 3033
rect 586 3003 589 3086
rect 602 3013 605 3093
rect 658 3046 661 3103
rect 658 3043 669 3046
rect 674 3043 677 3206
rect 714 3203 725 3206
rect 730 3203 733 3233
rect 1458 3226 1461 3246
rect 1786 3243 1797 3246
rect 762 3213 781 3216
rect 738 3203 749 3206
rect 690 3113 693 3136
rect 738 3123 741 3203
rect 762 3146 765 3196
rect 778 3146 781 3156
rect 762 3143 781 3146
rect 786 3133 789 3146
rect 778 3103 781 3126
rect 802 3123 805 3216
rect 818 3193 821 3206
rect 874 3183 877 3206
rect 922 3166 925 3216
rect 954 3193 957 3216
rect 818 3113 821 3136
rect 866 3123 869 3146
rect 898 3076 901 3126
rect 906 3123 909 3136
rect 914 3133 917 3166
rect 922 3163 949 3166
rect 946 3133 949 3163
rect 954 3143 957 3156
rect 970 3146 973 3216
rect 986 3203 989 3226
rect 1018 3183 1021 3206
rect 962 3133 965 3146
rect 970 3143 1013 3146
rect 970 3123 973 3143
rect 978 3133 989 3136
rect 890 3073 901 3076
rect 802 3053 829 3056
rect 610 3023 621 3026
rect 626 3023 653 3026
rect 650 3016 653 3023
rect 594 2996 597 3006
rect 586 2993 597 2996
rect 586 2903 589 2993
rect 594 2913 597 2986
rect 618 2946 621 2976
rect 626 2956 629 3006
rect 626 2953 637 2956
rect 618 2943 629 2946
rect 602 2933 621 2936
rect 626 2933 629 2943
rect 618 2926 621 2933
rect 610 2843 613 2926
rect 618 2923 629 2926
rect 634 2923 637 2946
rect 642 2926 645 3016
rect 650 3013 661 3016
rect 658 3003 661 3013
rect 642 2923 653 2926
rect 626 2903 629 2916
rect 650 2906 653 2923
rect 642 2903 653 2906
rect 546 2796 549 2806
rect 554 2803 565 2806
rect 570 2796 573 2806
rect 546 2793 573 2796
rect 570 2783 573 2793
rect 538 2753 573 2756
rect 498 2743 565 2746
rect 490 2733 517 2736
rect 514 2723 517 2733
rect 490 2686 493 2716
rect 522 2706 525 2736
rect 530 2733 549 2736
rect 554 2733 565 2736
rect 546 2726 549 2733
rect 538 2713 541 2726
rect 546 2723 557 2726
rect 514 2703 525 2706
rect 554 2703 557 2716
rect 490 2683 501 2686
rect 498 2616 501 2683
rect 490 2613 501 2616
rect 514 2616 517 2703
rect 562 2693 565 2733
rect 514 2613 525 2616
rect 490 2583 493 2613
rect 482 2553 493 2556
rect 418 2533 421 2546
rect 442 2543 453 2546
rect 450 2496 453 2543
rect 466 2523 469 2546
rect 386 2463 397 2466
rect 446 2493 453 2496
rect 386 2383 389 2463
rect 446 2446 449 2493
rect 434 2413 437 2446
rect 442 2443 449 2446
rect 378 2373 389 2376
rect 314 2363 341 2366
rect 282 2323 285 2363
rect 306 2323 309 2336
rect 210 2193 269 2196
rect 274 2186 277 2216
rect 210 2123 213 2186
rect 222 2183 277 2186
rect 282 2183 285 2206
rect 222 2116 225 2183
rect 234 2123 237 2136
rect 218 2113 225 2116
rect 162 1903 165 1916
rect 170 1813 173 1896
rect 146 1723 157 1726
rect 146 1683 149 1716
rect 154 1703 157 1723
rect 162 1716 165 1806
rect 170 1793 173 1806
rect 178 1776 181 1926
rect 186 1893 189 1926
rect 194 1923 205 1926
rect 194 1816 197 1923
rect 202 1903 205 1916
rect 186 1813 197 1816
rect 186 1783 189 1813
rect 178 1773 189 1776
rect 178 1723 181 1746
rect 186 1733 189 1773
rect 194 1733 197 1806
rect 202 1733 205 1826
rect 162 1713 173 1716
rect 154 1693 165 1696
rect 146 1613 149 1636
rect 154 1556 157 1676
rect 130 1553 157 1556
rect 130 1503 133 1553
rect 162 1546 165 1686
rect 170 1613 173 1713
rect 178 1563 181 1626
rect 146 1533 149 1546
rect 154 1543 165 1546
rect 138 1486 141 1526
rect 154 1523 157 1543
rect 170 1533 173 1556
rect 114 1106 117 1386
rect 122 1323 125 1396
rect 122 1303 125 1316
rect 122 1213 125 1226
rect 122 1173 125 1206
rect 122 1143 125 1166
rect 122 1113 125 1136
rect 114 1103 121 1106
rect 118 1036 121 1103
rect 118 1033 125 1036
rect 114 1003 117 1016
rect 106 923 117 926
rect 106 903 109 916
rect 114 896 117 923
rect 106 893 117 896
rect 106 783 109 893
rect 70 546 73 683
rect 70 543 77 546
rect 66 333 69 526
rect 74 513 77 543
rect 82 276 85 753
rect 90 716 93 736
rect 114 733 117 836
rect 98 723 109 726
rect 90 713 101 716
rect 90 603 93 696
rect 98 596 101 713
rect 114 706 117 726
rect 110 703 117 706
rect 110 646 113 703
rect 90 593 101 596
rect 106 643 113 646
rect 90 533 93 593
rect 106 493 109 643
rect 114 623 117 636
rect 122 523 125 1033
rect 130 1013 133 1486
rect 138 1483 157 1486
rect 138 1316 141 1476
rect 146 1413 149 1436
rect 146 1363 149 1406
rect 154 1356 157 1483
rect 162 1363 165 1426
rect 146 1353 157 1356
rect 146 1323 149 1353
rect 170 1346 173 1526
rect 178 1513 181 1526
rect 186 1503 189 1726
rect 194 1713 197 1726
rect 202 1626 205 1726
rect 194 1623 205 1626
rect 194 1613 197 1623
rect 194 1593 197 1606
rect 194 1496 197 1586
rect 178 1493 197 1496
rect 178 1403 181 1493
rect 170 1343 181 1346
rect 154 1333 165 1336
rect 138 1313 153 1316
rect 138 1253 141 1306
rect 150 1236 153 1313
rect 162 1303 165 1326
rect 170 1296 173 1336
rect 178 1323 181 1343
rect 162 1293 173 1296
rect 150 1233 157 1236
rect 138 1213 149 1216
rect 138 1203 149 1206
rect 146 1143 149 1156
rect 138 1073 141 1126
rect 146 1056 149 1136
rect 142 1053 149 1056
rect 130 933 133 946
rect 130 833 133 916
rect 142 846 145 1053
rect 142 843 149 846
rect 130 773 133 806
rect 130 693 133 756
rect 138 703 141 826
rect 138 683 141 696
rect 130 603 133 656
rect 130 533 133 546
rect 90 413 93 426
rect 98 403 101 416
rect 106 336 109 416
rect 122 413 125 516
rect 106 333 117 336
rect 122 333 125 346
rect 114 326 117 333
rect 106 313 109 326
rect 114 323 125 326
rect 130 323 133 336
rect 122 313 125 323
rect 130 296 133 316
rect 74 273 85 276
rect 122 293 133 296
rect 74 146 77 273
rect 90 156 93 266
rect 122 226 125 293
rect 98 213 101 226
rect 106 223 125 226
rect 106 203 109 223
rect 90 153 97 156
rect 74 143 85 146
rect 82 123 85 143
rect 94 106 97 153
rect 114 133 117 216
rect 138 123 141 646
rect 146 513 149 843
rect 154 623 157 1233
rect 162 1213 165 1293
rect 186 1266 189 1446
rect 194 1353 197 1486
rect 202 1453 205 1616
rect 202 1336 205 1416
rect 178 1263 189 1266
rect 198 1333 205 1336
rect 210 1333 213 2026
rect 218 2003 221 2113
rect 226 1973 229 2076
rect 242 2036 245 2156
rect 290 2153 293 2226
rect 338 2213 341 2363
rect 354 2216 357 2326
rect 386 2323 389 2373
rect 410 2323 413 2336
rect 442 2296 445 2443
rect 426 2293 445 2296
rect 354 2213 365 2216
rect 258 2106 261 2126
rect 266 2113 269 2136
rect 314 2133 325 2136
rect 258 2103 269 2106
rect 274 2103 277 2126
rect 290 2066 293 2116
rect 282 2063 293 2066
rect 238 2033 245 2036
rect 238 1976 241 2033
rect 250 2013 253 2026
rect 258 2003 261 2036
rect 282 2023 285 2063
rect 266 2013 285 2016
rect 238 1973 245 1976
rect 218 1953 237 1956
rect 242 1953 245 1973
rect 218 1933 221 1953
rect 250 1946 253 1996
rect 242 1943 253 1946
rect 218 1903 221 1916
rect 218 1803 221 1876
rect 226 1836 229 1936
rect 234 1893 237 1926
rect 242 1843 245 1943
rect 250 1933 261 1936
rect 250 1846 253 1933
rect 258 1913 261 1926
rect 266 1923 269 1956
rect 274 1896 277 2013
rect 282 1993 285 2006
rect 298 2003 301 2126
rect 306 2106 309 2126
rect 306 2103 313 2106
rect 310 1996 313 2103
rect 322 2096 325 2133
rect 330 2103 333 2206
rect 338 2193 341 2206
rect 362 2203 365 2213
rect 370 2156 373 2216
rect 354 2153 373 2156
rect 338 2096 341 2136
rect 322 2093 341 2096
rect 322 2016 325 2093
rect 338 2023 341 2056
rect 322 2013 341 2016
rect 346 2013 349 2126
rect 306 1993 313 1996
rect 322 2003 333 2006
rect 298 1933 301 1946
rect 306 1926 309 1993
rect 314 1933 317 1956
rect 282 1913 285 1926
rect 290 1903 293 1926
rect 298 1923 309 1926
rect 274 1893 281 1896
rect 250 1843 261 1846
rect 226 1833 253 1836
rect 226 1793 229 1816
rect 234 1763 237 1833
rect 258 1826 261 1843
rect 266 1833 269 1876
rect 278 1836 281 1893
rect 278 1833 285 1836
rect 242 1813 245 1826
rect 250 1823 261 1826
rect 218 1613 221 1736
rect 234 1733 237 1746
rect 242 1733 245 1806
rect 250 1743 253 1823
rect 258 1806 261 1816
rect 274 1813 277 1826
rect 258 1803 277 1806
rect 226 1623 229 1726
rect 218 1573 221 1606
rect 226 1593 229 1606
rect 218 1513 221 1536
rect 226 1523 229 1566
rect 218 1413 221 1506
rect 226 1413 229 1436
rect 226 1393 229 1406
rect 170 1233 173 1256
rect 162 953 165 1186
rect 170 1123 173 1226
rect 178 1116 181 1263
rect 198 1226 201 1333
rect 174 1113 181 1116
rect 186 1223 201 1226
rect 174 1036 177 1113
rect 170 1033 177 1036
rect 162 713 165 926
rect 170 813 173 1033
rect 178 873 181 1016
rect 186 913 189 1223
rect 210 1216 213 1326
rect 218 1276 221 1326
rect 226 1283 229 1326
rect 234 1323 237 1706
rect 242 1633 245 1726
rect 250 1623 253 1696
rect 258 1616 261 1726
rect 242 1533 245 1616
rect 250 1613 261 1616
rect 250 1533 253 1613
rect 242 1506 245 1526
rect 250 1513 253 1526
rect 242 1503 253 1506
rect 218 1273 237 1276
rect 202 1213 213 1216
rect 218 1213 221 1236
rect 194 1143 197 1156
rect 202 1143 205 1213
rect 210 1146 213 1206
rect 226 1203 229 1226
rect 234 1213 237 1273
rect 242 1243 245 1496
rect 250 1473 253 1503
rect 250 1233 253 1426
rect 242 1223 253 1226
rect 210 1143 229 1146
rect 202 1116 205 1136
rect 198 1113 205 1116
rect 198 1026 201 1113
rect 198 1023 205 1026
rect 194 993 197 1006
rect 194 893 197 936
rect 178 803 181 836
rect 186 823 197 826
rect 178 756 181 786
rect 170 753 181 756
rect 186 743 189 796
rect 194 783 197 816
rect 178 716 181 736
rect 170 713 181 716
rect 162 616 165 706
rect 170 686 173 706
rect 178 693 181 706
rect 170 683 177 686
rect 154 613 165 616
rect 162 413 165 556
rect 174 546 177 683
rect 186 653 189 716
rect 174 543 181 546
rect 178 416 181 543
rect 186 513 189 616
rect 194 433 197 716
rect 174 413 181 416
rect 146 323 149 386
rect 154 316 157 366
rect 146 313 157 316
rect 146 223 149 313
rect 162 233 165 336
rect 174 286 177 413
rect 186 296 189 406
rect 194 333 197 416
rect 202 393 205 1023
rect 210 1013 213 1136
rect 226 1123 229 1143
rect 234 1133 237 1146
rect 210 993 213 1006
rect 218 1003 221 1016
rect 210 866 213 926
rect 218 913 221 926
rect 226 916 229 1056
rect 234 923 237 1126
rect 226 913 237 916
rect 226 893 229 906
rect 234 903 237 913
rect 210 863 221 866
rect 210 813 213 826
rect 210 733 213 806
rect 218 733 221 863
rect 210 703 213 726
rect 218 693 221 706
rect 226 656 229 816
rect 234 793 237 886
rect 242 803 245 1223
rect 250 1193 253 1216
rect 258 1163 261 1606
rect 266 1523 269 1736
rect 274 1583 277 1803
rect 282 1713 285 1833
rect 274 1523 277 1546
rect 266 1483 269 1516
rect 266 1386 269 1466
rect 274 1433 277 1446
rect 274 1396 277 1426
rect 282 1403 285 1706
rect 290 1686 293 1846
rect 298 1723 301 1923
rect 314 1903 317 1926
rect 322 1896 325 2003
rect 338 1966 341 2013
rect 354 2003 357 2153
rect 378 2136 381 2226
rect 386 2143 389 2166
rect 370 2133 381 2136
rect 394 2133 397 2246
rect 362 1996 365 2106
rect 306 1893 325 1896
rect 330 1963 341 1966
rect 354 1993 365 1996
rect 306 1733 309 1893
rect 322 1833 325 1876
rect 330 1826 333 1963
rect 338 1843 341 1936
rect 346 1913 349 1926
rect 314 1823 333 1826
rect 314 1813 317 1823
rect 338 1813 341 1826
rect 322 1726 325 1736
rect 330 1733 333 1776
rect 338 1733 341 1806
rect 346 1793 349 1906
rect 306 1723 325 1726
rect 306 1703 309 1723
rect 322 1703 325 1716
rect 290 1683 321 1686
rect 290 1603 293 1646
rect 306 1613 309 1676
rect 318 1626 321 1683
rect 318 1623 325 1626
rect 298 1603 309 1606
rect 290 1413 293 1566
rect 298 1423 301 1603
rect 306 1543 309 1586
rect 314 1533 317 1606
rect 322 1546 325 1623
rect 330 1613 333 1726
rect 338 1713 341 1726
rect 330 1553 333 1586
rect 338 1556 341 1706
rect 346 1563 349 1616
rect 354 1606 357 1993
rect 370 1946 373 2133
rect 378 2033 381 2126
rect 386 2113 389 2126
rect 402 2043 405 2216
rect 418 2183 421 2206
rect 418 2126 421 2136
rect 410 2123 421 2126
rect 426 2123 429 2293
rect 410 2023 413 2123
rect 418 2073 421 2116
rect 378 1983 381 2016
rect 394 2003 397 2016
rect 386 1973 389 1996
rect 402 1946 405 2016
rect 410 1963 413 2006
rect 362 1943 373 1946
rect 394 1943 405 1946
rect 362 1896 365 1943
rect 370 1933 389 1936
rect 370 1923 381 1926
rect 378 1903 381 1923
rect 362 1893 373 1896
rect 362 1823 365 1886
rect 362 1713 365 1816
rect 362 1613 365 1626
rect 354 1603 365 1606
rect 338 1553 349 1556
rect 322 1543 341 1546
rect 306 1463 309 1526
rect 274 1393 293 1396
rect 306 1393 309 1416
rect 314 1403 317 1526
rect 322 1513 325 1526
rect 330 1523 333 1536
rect 322 1436 325 1506
rect 330 1443 333 1466
rect 322 1433 333 1436
rect 322 1413 325 1426
rect 330 1396 333 1433
rect 314 1393 333 1396
rect 266 1383 277 1386
rect 250 923 253 1126
rect 258 1053 261 1156
rect 266 1123 269 1356
rect 274 1133 277 1383
rect 282 1323 285 1386
rect 290 1353 293 1393
rect 290 1333 293 1346
rect 298 1333 301 1376
rect 282 1303 285 1316
rect 290 1246 293 1326
rect 282 1243 293 1246
rect 282 1116 285 1243
rect 290 1176 293 1236
rect 298 1226 301 1326
rect 306 1303 309 1326
rect 306 1233 309 1266
rect 298 1223 309 1226
rect 298 1193 301 1216
rect 290 1173 297 1176
rect 278 1113 285 1116
rect 250 833 253 916
rect 258 913 261 1026
rect 266 913 269 1046
rect 278 1036 281 1113
rect 294 1106 297 1173
rect 306 1133 309 1223
rect 314 1213 317 1393
rect 322 1263 325 1356
rect 330 1333 333 1386
rect 322 1233 325 1246
rect 314 1183 317 1206
rect 330 1196 333 1326
rect 322 1193 333 1196
rect 322 1173 325 1193
rect 290 1103 297 1106
rect 278 1033 285 1036
rect 258 863 261 906
rect 258 786 261 856
rect 266 813 269 876
rect 266 793 269 806
rect 210 653 229 656
rect 210 606 213 653
rect 234 646 237 786
rect 258 783 269 786
rect 250 726 253 776
rect 242 723 253 726
rect 218 643 237 646
rect 218 613 221 643
rect 226 613 237 616
rect 210 603 221 606
rect 218 556 221 603
rect 226 593 229 606
rect 242 586 245 696
rect 258 666 261 726
rect 234 583 245 586
rect 250 663 261 666
rect 218 553 225 556
rect 210 523 213 546
rect 210 413 213 516
rect 222 476 225 553
rect 218 473 225 476
rect 194 303 197 316
rect 210 313 213 356
rect 186 293 205 296
rect 174 283 181 286
rect 170 213 173 246
rect 178 223 181 283
rect 178 203 181 216
rect 194 203 197 216
rect 186 133 189 196
rect 202 133 205 293
rect 210 133 213 226
rect 218 216 221 473
rect 234 456 237 583
rect 250 506 253 663
rect 258 523 261 656
rect 266 516 269 783
rect 274 633 277 1016
rect 282 853 285 1033
rect 290 1023 293 1103
rect 306 1023 309 1126
rect 322 1113 325 1136
rect 330 1123 333 1186
rect 338 1173 341 1543
rect 346 1413 349 1553
rect 354 1443 357 1576
rect 346 1393 349 1406
rect 354 1403 357 1416
rect 346 1366 349 1386
rect 362 1373 365 1603
rect 370 1533 373 1893
rect 378 1833 381 1856
rect 378 1723 381 1826
rect 386 1823 389 1933
rect 386 1733 389 1796
rect 394 1776 397 1943
rect 402 1923 405 1936
rect 402 1913 413 1916
rect 418 1913 421 2056
rect 426 2003 429 2096
rect 434 2013 437 2286
rect 442 2116 445 2226
rect 450 2203 453 2326
rect 458 2323 461 2406
rect 490 2386 493 2553
rect 498 2543 509 2546
rect 506 2533 509 2543
rect 506 2493 509 2526
rect 514 2503 517 2596
rect 522 2516 525 2613
rect 530 2573 533 2686
rect 538 2523 541 2616
rect 522 2513 541 2516
rect 482 2383 493 2386
rect 482 2296 485 2383
rect 498 2306 501 2416
rect 538 2413 541 2513
rect 546 2506 549 2656
rect 570 2646 573 2753
rect 578 2653 581 2826
rect 594 2796 597 2816
rect 590 2793 597 2796
rect 590 2696 593 2793
rect 618 2766 621 2856
rect 602 2763 621 2766
rect 602 2703 605 2763
rect 590 2693 597 2696
rect 570 2643 581 2646
rect 554 2603 557 2626
rect 562 2606 565 2626
rect 570 2613 573 2636
rect 562 2603 573 2606
rect 578 2596 581 2643
rect 586 2603 589 2616
rect 562 2583 565 2596
rect 578 2593 589 2596
rect 546 2503 557 2506
rect 506 2323 509 2386
rect 522 2323 525 2336
rect 498 2303 505 2306
rect 482 2293 493 2296
rect 458 2183 461 2256
rect 450 2133 469 2136
rect 474 2133 477 2146
rect 482 2143 485 2156
rect 466 2126 469 2133
rect 442 2113 449 2116
rect 446 2006 449 2113
rect 458 2083 461 2126
rect 466 2123 477 2126
rect 474 2103 477 2116
rect 482 2096 485 2126
rect 490 2113 493 2293
rect 502 2216 505 2303
rect 502 2213 509 2216
rect 506 2203 509 2213
rect 498 2123 501 2176
rect 482 2093 489 2096
rect 442 2003 449 2006
rect 442 1933 445 2003
rect 458 1983 461 1996
rect 466 1953 469 2016
rect 474 1946 477 2056
rect 486 2036 489 2093
rect 506 2066 509 2136
rect 498 2063 509 2066
rect 486 2033 493 2036
rect 482 2003 485 2026
rect 450 1943 477 1946
rect 410 1906 413 1913
rect 410 1903 429 1906
rect 402 1783 405 1896
rect 410 1813 413 1826
rect 394 1773 405 1776
rect 378 1643 381 1716
rect 402 1646 405 1773
rect 418 1713 421 1876
rect 434 1823 437 1926
rect 442 1853 445 1926
rect 450 1923 453 1943
rect 458 1916 461 1936
rect 482 1933 485 1966
rect 490 1933 493 2033
rect 454 1913 461 1916
rect 474 1913 477 1926
rect 454 1826 457 1913
rect 426 1793 429 1816
rect 442 1813 445 1826
rect 450 1823 457 1826
rect 434 1803 445 1806
rect 426 1723 429 1736
rect 434 1733 437 1803
rect 450 1796 453 1823
rect 466 1813 469 1906
rect 482 1876 485 1896
rect 478 1873 485 1876
rect 442 1793 453 1796
rect 442 1716 445 1793
rect 450 1733 453 1746
rect 398 1643 405 1646
rect 378 1613 381 1636
rect 378 1593 381 1606
rect 386 1603 389 1626
rect 386 1533 389 1576
rect 398 1566 401 1643
rect 426 1636 429 1716
rect 410 1633 429 1636
rect 438 1713 445 1716
rect 398 1563 405 1566
rect 370 1523 381 1526
rect 386 1473 389 1526
rect 370 1463 389 1466
rect 370 1443 373 1463
rect 370 1413 373 1426
rect 378 1423 381 1456
rect 386 1443 389 1463
rect 378 1413 389 1416
rect 346 1363 353 1366
rect 350 1236 353 1363
rect 362 1313 365 1346
rect 346 1233 353 1236
rect 338 1033 341 1166
rect 346 1153 349 1233
rect 354 1203 357 1216
rect 362 1186 365 1266
rect 370 1203 373 1406
rect 378 1343 381 1413
rect 378 1186 381 1336
rect 386 1333 389 1406
rect 386 1203 389 1326
rect 354 1183 365 1186
rect 370 1183 381 1186
rect 346 1123 349 1136
rect 354 1103 357 1183
rect 386 1176 389 1196
rect 314 1023 349 1026
rect 314 1016 317 1023
rect 354 1016 357 1066
rect 298 1013 317 1016
rect 290 966 293 1006
rect 290 963 301 966
rect 282 813 285 846
rect 282 733 285 806
rect 290 733 293 956
rect 298 826 301 963
rect 306 923 309 936
rect 306 843 309 916
rect 314 873 317 1013
rect 322 1003 325 1016
rect 330 946 333 1006
rect 338 953 341 1016
rect 346 1013 357 1016
rect 346 946 349 1013
rect 362 996 365 1176
rect 330 943 349 946
rect 358 993 365 996
rect 370 1173 389 1176
rect 358 936 361 993
rect 330 933 361 936
rect 298 823 317 826
rect 298 783 301 816
rect 274 603 277 626
rect 226 453 237 456
rect 246 503 253 506
rect 258 513 269 516
rect 274 516 277 576
rect 282 533 285 706
rect 290 646 293 706
rect 298 693 301 776
rect 306 653 309 816
rect 314 746 317 823
rect 322 803 325 916
rect 330 863 333 926
rect 338 843 341 926
rect 330 833 341 836
rect 330 773 333 826
rect 314 743 333 746
rect 314 703 317 736
rect 322 703 325 716
rect 330 686 333 743
rect 326 683 333 686
rect 290 643 317 646
rect 290 603 293 643
rect 306 623 309 636
rect 298 543 301 616
rect 306 553 309 616
rect 314 603 317 643
rect 326 626 329 683
rect 322 623 329 626
rect 274 513 285 516
rect 226 333 229 453
rect 234 403 237 436
rect 246 426 249 503
rect 242 423 249 426
rect 242 386 245 423
rect 238 383 245 386
rect 226 233 229 326
rect 238 266 241 383
rect 250 363 253 416
rect 258 403 261 513
rect 258 356 261 396
rect 250 353 261 356
rect 238 263 245 266
rect 242 243 245 263
rect 218 213 229 216
rect 226 166 229 213
rect 218 163 229 166
rect 218 126 221 163
rect 186 123 197 126
rect 210 123 221 126
rect 186 116 189 123
rect 170 113 189 116
rect 250 113 253 353
rect 266 326 269 506
rect 282 376 285 513
rect 298 493 301 536
rect 314 533 317 566
rect 322 546 325 623
rect 330 603 333 616
rect 322 543 333 546
rect 306 513 309 526
rect 314 496 317 526
rect 322 513 325 536
rect 330 506 333 543
rect 338 523 341 833
rect 346 623 349 926
rect 354 916 357 933
rect 354 913 361 916
rect 358 856 361 913
rect 354 853 361 856
rect 354 793 357 853
rect 362 803 365 836
rect 354 733 357 786
rect 370 736 373 1173
rect 378 893 381 1136
rect 386 1133 389 1166
rect 386 1113 389 1126
rect 386 1006 389 1106
rect 394 1083 397 1546
rect 402 1323 405 1563
rect 410 1413 413 1633
rect 418 1623 429 1626
rect 418 1523 421 1623
rect 438 1616 441 1713
rect 426 1613 441 1616
rect 418 1503 421 1516
rect 418 1423 421 1446
rect 418 1393 421 1406
rect 426 1396 429 1613
rect 434 1543 437 1606
rect 450 1536 453 1726
rect 458 1723 461 1806
rect 466 1753 469 1806
rect 478 1756 481 1873
rect 490 1846 493 1926
rect 498 1913 501 2063
rect 506 2013 509 2056
rect 514 1966 517 2236
rect 522 2143 525 2226
rect 530 2203 533 2216
rect 538 2166 541 2296
rect 546 2216 549 2326
rect 554 2293 557 2503
rect 562 2483 565 2556
rect 586 2516 589 2593
rect 594 2523 597 2693
rect 610 2636 613 2756
rect 618 2733 621 2746
rect 626 2663 629 2866
rect 642 2846 645 2903
rect 658 2853 661 2966
rect 666 2956 669 3043
rect 802 3036 805 3053
rect 674 3013 677 3026
rect 682 2993 685 3016
rect 698 3013 701 3036
rect 706 3033 805 3036
rect 690 2973 693 3006
rect 706 3003 709 3033
rect 714 2966 717 3016
rect 722 3003 725 3016
rect 738 3013 741 3026
rect 730 2973 733 3006
rect 746 3003 749 3033
rect 698 2963 741 2966
rect 666 2953 677 2956
rect 674 2866 677 2953
rect 698 2923 701 2963
rect 666 2863 677 2866
rect 666 2846 669 2863
rect 642 2843 653 2846
rect 650 2823 653 2843
rect 658 2843 669 2846
rect 658 2813 661 2843
rect 666 2813 669 2836
rect 634 2743 637 2806
rect 674 2803 677 2846
rect 706 2836 709 2946
rect 698 2833 709 2836
rect 682 2813 709 2816
rect 714 2813 717 2936
rect 722 2933 733 2936
rect 722 2886 725 2926
rect 730 2903 733 2933
rect 738 2923 741 2963
rect 754 2926 757 3016
rect 778 3013 781 3026
rect 762 2973 765 3006
rect 794 2983 797 3016
rect 802 3003 805 3033
rect 810 2946 813 3046
rect 826 3006 829 3053
rect 842 3013 845 3056
rect 890 3026 893 3073
rect 882 3023 893 3026
rect 850 3013 861 3016
rect 826 3003 869 3006
rect 834 2976 837 2996
rect 794 2943 813 2946
rect 826 2973 837 2976
rect 762 2933 773 2936
rect 794 2926 797 2943
rect 802 2933 821 2936
rect 826 2933 829 2973
rect 834 2933 837 2956
rect 866 2953 869 3003
rect 874 2983 877 3006
rect 882 2946 885 3023
rect 898 2993 901 3016
rect 850 2943 885 2946
rect 818 2926 821 2933
rect 746 2923 765 2926
rect 746 2916 749 2923
rect 778 2916 781 2926
rect 794 2923 813 2926
rect 818 2923 845 2926
rect 738 2913 749 2916
rect 754 2913 781 2916
rect 722 2883 729 2886
rect 690 2746 693 2806
rect 650 2743 693 2746
rect 634 2713 637 2736
rect 650 2733 653 2743
rect 658 2733 669 2736
rect 610 2633 617 2636
rect 602 2613 605 2626
rect 602 2553 605 2606
rect 614 2576 617 2633
rect 642 2626 645 2726
rect 658 2646 661 2726
rect 674 2723 677 2736
rect 690 2733 693 2743
rect 698 2733 701 2766
rect 626 2603 629 2626
rect 634 2623 645 2626
rect 654 2643 661 2646
rect 610 2573 617 2576
rect 602 2523 605 2546
rect 586 2513 597 2516
rect 594 2466 597 2513
rect 594 2463 605 2466
rect 578 2366 581 2406
rect 570 2363 581 2366
rect 570 2323 573 2363
rect 602 2323 605 2463
rect 554 2223 557 2236
rect 570 2233 597 2236
rect 546 2213 557 2216
rect 554 2203 557 2213
rect 562 2203 565 2216
rect 570 2213 573 2233
rect 578 2223 589 2226
rect 534 2163 541 2166
rect 522 2073 525 2126
rect 522 2023 525 2066
rect 534 2046 537 2163
rect 546 2133 549 2156
rect 534 2043 541 2046
rect 530 2003 533 2026
rect 538 2023 541 2043
rect 514 1963 525 1966
rect 490 1843 501 1846
rect 478 1753 485 1756
rect 474 1726 477 1736
rect 482 1733 485 1753
rect 466 1723 477 1726
rect 458 1653 461 1716
rect 434 1533 453 1536
rect 434 1453 437 1516
rect 442 1463 445 1526
rect 450 1473 453 1516
rect 442 1413 445 1446
rect 450 1413 453 1456
rect 434 1403 453 1406
rect 426 1393 437 1396
rect 410 1333 429 1336
rect 434 1333 437 1393
rect 402 1293 405 1316
rect 402 1203 405 1246
rect 402 1093 405 1176
rect 394 1013 405 1016
rect 386 1003 397 1006
rect 386 916 389 996
rect 394 923 397 1003
rect 402 933 405 1013
rect 410 986 413 1316
rect 418 1123 421 1296
rect 418 1003 421 1096
rect 426 1003 429 1333
rect 434 1296 437 1326
rect 442 1303 445 1366
rect 434 1293 445 1296
rect 434 1123 437 1256
rect 442 1243 445 1293
rect 450 1236 453 1403
rect 442 1233 453 1236
rect 442 1153 445 1233
rect 450 1213 453 1226
rect 442 1113 445 1136
rect 450 1103 453 1206
rect 458 1096 461 1606
rect 466 1383 469 1723
rect 474 1603 477 1716
rect 474 1506 477 1566
rect 482 1513 485 1666
rect 474 1503 485 1506
rect 466 1293 469 1336
rect 466 1233 469 1286
rect 474 1226 477 1476
rect 482 1453 485 1503
rect 482 1403 485 1446
rect 482 1363 485 1396
rect 490 1383 493 1826
rect 498 1803 501 1843
rect 498 1773 501 1796
rect 498 1613 501 1766
rect 498 1593 501 1606
rect 498 1543 501 1576
rect 498 1356 501 1536
rect 466 1223 477 1226
rect 482 1353 501 1356
rect 466 1146 469 1223
rect 474 1196 477 1216
rect 482 1203 485 1353
rect 474 1193 485 1196
rect 466 1143 477 1146
rect 434 1006 437 1096
rect 442 1093 461 1096
rect 442 1013 445 1093
rect 434 1003 441 1006
rect 410 983 417 986
rect 386 913 405 916
rect 378 793 381 816
rect 366 733 373 736
rect 310 493 317 496
rect 322 503 333 506
rect 310 426 313 493
rect 310 423 317 426
rect 258 323 269 326
rect 274 373 285 376
rect 258 223 261 323
rect 274 316 277 373
rect 298 356 301 416
rect 306 393 309 406
rect 282 353 301 356
rect 266 313 277 316
rect 298 316 301 326
rect 314 323 317 423
rect 322 333 325 503
rect 322 316 325 326
rect 298 313 325 316
rect 266 216 269 313
rect 330 306 333 426
rect 314 286 317 306
rect 306 283 317 286
rect 322 303 333 306
rect 338 303 341 496
rect 346 313 349 596
rect 354 353 357 726
rect 366 676 369 733
rect 378 713 381 726
rect 378 686 381 706
rect 386 696 389 913
rect 414 906 417 983
rect 438 946 441 1003
rect 438 943 445 946
rect 410 903 417 906
rect 426 903 429 936
rect 434 913 437 926
rect 394 706 397 846
rect 402 803 405 826
rect 410 773 413 903
rect 402 723 413 726
rect 402 713 405 723
rect 394 703 405 706
rect 386 693 397 696
rect 378 683 389 686
rect 366 673 373 676
rect 362 433 365 656
rect 370 523 373 673
rect 378 463 381 606
rect 386 596 389 656
rect 394 603 397 693
rect 402 643 405 703
rect 418 656 421 886
rect 426 723 429 896
rect 442 893 445 943
rect 434 863 445 866
rect 434 813 437 863
rect 434 783 437 806
rect 442 793 445 816
rect 434 716 437 776
rect 410 653 421 656
rect 426 713 437 716
rect 386 593 397 596
rect 378 426 381 436
rect 362 423 381 426
rect 362 413 365 423
rect 370 413 381 416
rect 362 303 365 406
rect 378 396 381 413
rect 374 393 381 396
rect 374 316 377 393
rect 386 323 389 526
rect 394 386 397 593
rect 402 513 405 616
rect 410 603 413 653
rect 418 583 421 646
rect 426 576 429 713
rect 434 623 437 676
rect 422 573 429 576
rect 410 533 413 546
rect 422 526 425 573
rect 418 523 425 526
rect 402 413 405 436
rect 418 413 421 523
rect 434 506 437 606
rect 442 586 445 736
rect 450 603 453 1086
rect 466 1053 469 1136
rect 458 1016 461 1036
rect 458 1013 469 1016
rect 458 923 461 1006
rect 458 633 461 916
rect 466 723 469 946
rect 466 633 469 696
rect 474 653 477 1143
rect 482 1093 485 1193
rect 482 1013 485 1076
rect 482 813 485 1006
rect 490 936 493 1336
rect 506 1333 509 1936
rect 514 1933 517 1956
rect 514 1913 517 1926
rect 522 1906 525 1963
rect 530 1923 533 1936
rect 514 1603 517 1906
rect 522 1903 529 1906
rect 526 1846 529 1903
rect 522 1843 529 1846
rect 522 1736 525 1843
rect 538 1826 541 2016
rect 546 1963 549 2126
rect 530 1823 541 1826
rect 530 1743 533 1823
rect 546 1816 549 1876
rect 554 1826 557 2146
rect 562 2143 565 2156
rect 570 2133 573 2176
rect 562 2093 565 2126
rect 562 1953 565 2046
rect 578 2036 581 2223
rect 586 2203 589 2216
rect 594 2196 597 2233
rect 602 2203 605 2316
rect 610 2196 613 2573
rect 634 2533 637 2623
rect 642 2583 645 2606
rect 654 2596 657 2643
rect 666 2623 669 2636
rect 666 2603 669 2616
rect 674 2613 677 2646
rect 682 2616 685 2726
rect 706 2643 709 2813
rect 714 2743 717 2806
rect 726 2776 729 2883
rect 738 2803 741 2896
rect 778 2893 781 2913
rect 746 2813 757 2816
rect 722 2773 729 2776
rect 722 2753 725 2773
rect 746 2766 749 2796
rect 754 2773 757 2806
rect 762 2783 765 2806
rect 746 2763 757 2766
rect 754 2733 757 2763
rect 770 2743 773 2826
rect 778 2796 781 2816
rect 778 2793 789 2796
rect 786 2746 789 2793
rect 778 2743 789 2746
rect 802 2746 805 2836
rect 810 2753 813 2923
rect 834 2896 837 2916
rect 842 2903 845 2923
rect 830 2893 837 2896
rect 818 2803 821 2866
rect 830 2826 833 2893
rect 830 2823 837 2826
rect 826 2783 829 2806
rect 802 2743 813 2746
rect 754 2713 757 2726
rect 762 2723 765 2736
rect 778 2706 781 2743
rect 770 2703 781 2706
rect 682 2613 701 2616
rect 714 2613 717 2626
rect 746 2623 749 2636
rect 654 2593 661 2596
rect 658 2536 661 2593
rect 674 2583 677 2606
rect 690 2603 701 2606
rect 706 2583 709 2606
rect 650 2533 661 2536
rect 690 2533 693 2576
rect 714 2533 717 2546
rect 722 2533 725 2556
rect 650 2516 653 2533
rect 646 2513 653 2516
rect 618 2396 621 2416
rect 618 2393 625 2396
rect 622 2316 625 2393
rect 646 2376 649 2513
rect 658 2413 661 2526
rect 666 2486 669 2506
rect 666 2483 677 2486
rect 674 2416 677 2483
rect 698 2446 701 2526
rect 730 2513 733 2616
rect 746 2536 749 2606
rect 754 2603 757 2666
rect 770 2586 773 2703
rect 786 2663 789 2726
rect 802 2713 805 2736
rect 778 2603 781 2616
rect 794 2603 797 2626
rect 802 2613 805 2646
rect 738 2533 749 2536
rect 762 2583 773 2586
rect 738 2513 741 2533
rect 762 2456 765 2583
rect 778 2553 781 2596
rect 810 2546 813 2743
rect 834 2736 837 2823
rect 826 2733 837 2736
rect 842 2733 845 2876
rect 850 2813 853 2943
rect 866 2933 885 2936
rect 890 2933 893 2976
rect 882 2926 885 2933
rect 858 2873 861 2926
rect 866 2903 869 2926
rect 882 2923 893 2926
rect 882 2913 893 2916
rect 890 2876 893 2913
rect 898 2893 901 2936
rect 890 2873 897 2876
rect 858 2733 861 2816
rect 866 2736 869 2816
rect 874 2763 877 2826
rect 882 2803 885 2866
rect 894 2816 897 2873
rect 894 2813 901 2816
rect 906 2813 909 3106
rect 914 2883 917 3116
rect 946 3113 957 3116
rect 922 3043 957 3046
rect 922 3003 925 3043
rect 930 2986 933 3016
rect 938 3003 941 3036
rect 946 3003 949 3016
rect 922 2983 933 2986
rect 922 2853 925 2983
rect 930 2896 933 2936
rect 938 2906 941 2926
rect 946 2913 949 2926
rect 954 2916 957 3043
rect 962 2983 965 3006
rect 978 3003 981 3126
rect 1002 3113 1005 3136
rect 1010 3123 1013 3143
rect 1018 3133 1021 3166
rect 1066 3133 1069 3216
rect 1098 3213 1101 3226
rect 1458 3223 1465 3226
rect 1122 3193 1125 3206
rect 1074 3133 1077 3156
rect 1106 3143 1109 3166
rect 1098 3126 1101 3136
rect 1018 3113 1021 3126
rect 1058 3123 1069 3126
rect 1090 3123 1101 3126
rect 1058 3106 1061 3123
rect 1090 3116 1093 3123
rect 1066 3113 1093 3116
rect 1058 3103 1069 3106
rect 1098 3103 1101 3116
rect 1042 3016 1045 3066
rect 986 2963 989 3016
rect 994 2933 997 3006
rect 1010 2953 1013 3016
rect 1042 3013 1049 3016
rect 1018 2946 1021 3006
rect 1026 3003 1037 3006
rect 1026 2983 1029 3003
rect 1034 2973 1037 2996
rect 1046 2966 1049 3013
rect 1058 2986 1061 3016
rect 1066 3003 1069 3103
rect 1106 3063 1109 3136
rect 1130 3123 1133 3216
rect 1154 3183 1157 3206
rect 1138 3133 1141 3176
rect 1186 3133 1189 3216
rect 1234 3193 1237 3216
rect 1258 3156 1261 3216
rect 1266 3203 1277 3206
rect 1290 3183 1293 3206
rect 1186 3113 1189 3126
rect 1194 3113 1197 3136
rect 1202 3076 1205 3126
rect 1218 3123 1221 3136
rect 1234 3133 1237 3146
rect 1218 3103 1221 3116
rect 1202 3073 1213 3076
rect 1074 3013 1077 3046
rect 1090 3023 1117 3026
rect 1090 3013 1093 3023
rect 1122 3013 1125 3056
rect 1130 3006 1133 3036
rect 1138 3016 1141 3026
rect 1138 3013 1157 3016
rect 1162 3013 1165 3036
rect 1082 2993 1085 3006
rect 1090 2986 1093 3006
rect 1130 3003 1149 3006
rect 1058 2983 1093 2986
rect 1074 2966 1077 2983
rect 1046 2963 1053 2966
rect 1018 2943 1037 2946
rect 1002 2933 1029 2936
rect 1002 2926 1005 2933
rect 970 2923 981 2926
rect 954 2913 965 2916
rect 938 2903 965 2906
rect 970 2903 973 2916
rect 930 2893 957 2896
rect 938 2813 941 2836
rect 866 2733 877 2736
rect 818 2713 821 2726
rect 826 2693 829 2733
rect 834 2723 845 2726
rect 818 2603 821 2616
rect 826 2613 829 2676
rect 826 2596 829 2606
rect 834 2603 837 2723
rect 842 2713 853 2716
rect 842 2613 845 2636
rect 850 2596 853 2626
rect 858 2613 861 2706
rect 866 2606 869 2726
rect 826 2593 853 2596
rect 858 2603 869 2606
rect 858 2583 861 2603
rect 874 2566 877 2733
rect 882 2686 885 2736
rect 890 2726 893 2806
rect 898 2756 901 2813
rect 930 2783 933 2806
rect 946 2773 949 2816
rect 898 2753 925 2756
rect 898 2733 909 2736
rect 914 2733 917 2746
rect 922 2726 925 2753
rect 938 2733 941 2746
rect 890 2723 901 2726
rect 890 2703 893 2716
rect 882 2683 889 2686
rect 886 2606 889 2683
rect 866 2563 877 2566
rect 882 2603 889 2606
rect 810 2543 821 2546
rect 786 2483 789 2536
rect 818 2496 821 2543
rect 834 2523 837 2546
rect 810 2493 821 2496
rect 866 2496 869 2563
rect 866 2493 877 2496
rect 762 2453 773 2456
rect 698 2443 709 2446
rect 666 2413 677 2416
rect 706 2413 709 2443
rect 666 2383 669 2413
rect 634 2373 649 2376
rect 714 2376 717 2406
rect 730 2403 733 2416
rect 754 2376 757 2416
rect 714 2373 757 2376
rect 634 2323 637 2373
rect 642 2333 653 2336
rect 642 2316 645 2333
rect 690 2323 693 2336
rect 622 2313 645 2316
rect 618 2213 621 2306
rect 650 2296 653 2316
rect 714 2313 717 2326
rect 650 2293 661 2296
rect 634 2213 637 2276
rect 658 2236 661 2293
rect 642 2206 645 2236
rect 626 2203 645 2206
rect 650 2233 661 2236
rect 650 2196 653 2233
rect 722 2216 725 2336
rect 594 2193 613 2196
rect 642 2193 653 2196
rect 594 2123 597 2136
rect 602 2123 605 2193
rect 586 2103 589 2116
rect 570 2033 581 2036
rect 570 1936 573 2033
rect 578 1946 581 2026
rect 586 2003 589 2026
rect 594 2003 597 2096
rect 602 2013 605 2116
rect 578 1943 589 1946
rect 562 1923 565 1936
rect 570 1933 581 1936
rect 562 1856 565 1916
rect 570 1893 573 1926
rect 578 1863 581 1933
rect 562 1853 573 1856
rect 554 1823 565 1826
rect 538 1803 541 1816
rect 546 1813 557 1816
rect 522 1733 533 1736
rect 522 1633 525 1726
rect 514 1523 517 1596
rect 514 1483 517 1516
rect 522 1463 525 1616
rect 530 1426 533 1733
rect 538 1723 541 1796
rect 546 1783 549 1806
rect 554 1743 557 1796
rect 562 1746 565 1823
rect 570 1756 573 1853
rect 578 1813 581 1846
rect 586 1793 589 1943
rect 594 1923 597 1956
rect 602 1923 605 1936
rect 610 1903 613 2146
rect 618 2016 621 2116
rect 626 2033 629 2136
rect 618 2013 625 2016
rect 622 1936 625 2013
rect 634 2003 637 2126
rect 642 1966 645 2193
rect 650 2043 653 2186
rect 658 2026 661 2216
rect 666 2163 669 2206
rect 666 2133 669 2156
rect 666 2026 669 2036
rect 650 1983 653 2026
rect 658 2023 669 2026
rect 674 2026 677 2216
rect 714 2213 725 2216
rect 682 2143 685 2206
rect 682 2093 685 2136
rect 690 2123 693 2186
rect 714 2166 717 2213
rect 738 2176 741 2206
rect 762 2196 765 2376
rect 770 2323 773 2453
rect 810 2353 813 2493
rect 874 2473 877 2493
rect 882 2456 885 2603
rect 898 2586 901 2723
rect 914 2713 917 2726
rect 922 2723 941 2726
rect 946 2723 949 2746
rect 954 2733 957 2893
rect 978 2836 981 2923
rect 994 2923 1005 2926
rect 1010 2923 1021 2926
rect 1034 2923 1037 2943
rect 994 2913 997 2923
rect 1050 2916 1053 2963
rect 1042 2913 1053 2916
rect 1066 2963 1077 2966
rect 970 2833 981 2836
rect 970 2776 973 2833
rect 986 2813 989 2826
rect 1002 2803 1005 2886
rect 1042 2813 1045 2913
rect 1066 2906 1069 2963
rect 1082 2916 1085 2936
rect 1090 2926 1093 2976
rect 1098 2933 1101 2946
rect 1106 2933 1109 2956
rect 1114 2953 1141 2956
rect 1114 2926 1117 2953
rect 1090 2923 1101 2926
rect 1106 2923 1117 2926
rect 1106 2916 1109 2923
rect 1082 2913 1109 2916
rect 1066 2903 1077 2906
rect 1074 2863 1077 2903
rect 1082 2813 1085 2826
rect 1090 2793 1093 2816
rect 1122 2813 1125 2946
rect 1138 2923 1141 2953
rect 1146 2853 1149 2996
rect 1154 2933 1157 3013
rect 1162 2983 1165 3006
rect 1210 3003 1213 3073
rect 1162 2943 1165 2966
rect 1218 2936 1221 3016
rect 1234 3013 1237 3056
rect 1226 2993 1229 3006
rect 1226 2943 1229 2966
rect 1234 2953 1237 3006
rect 1242 2996 1245 3146
rect 1250 3116 1253 3156
rect 1258 3153 1301 3156
rect 1266 3133 1269 3146
rect 1250 3113 1261 3116
rect 1258 3026 1261 3113
rect 1274 3063 1277 3126
rect 1250 3023 1261 3026
rect 1250 3003 1253 3023
rect 1242 2993 1253 2996
rect 1250 2973 1253 2993
rect 1266 2983 1269 3006
rect 1274 2946 1277 2966
rect 1282 2956 1285 3136
rect 1298 3123 1301 3153
rect 1306 3133 1309 3176
rect 1330 3133 1333 3216
rect 1370 3203 1373 3216
rect 1394 3183 1397 3206
rect 1386 3153 1421 3156
rect 1346 3133 1349 3146
rect 1370 3126 1373 3136
rect 1290 3013 1293 3046
rect 1282 2953 1293 2956
rect 1298 2953 1301 3026
rect 1306 3003 1309 3016
rect 1314 3003 1317 3016
rect 1330 3013 1333 3126
rect 1362 3123 1373 3126
rect 1362 3116 1365 3123
rect 1338 3113 1365 3116
rect 1370 3093 1373 3116
rect 1378 3113 1381 3136
rect 1386 3103 1389 3153
rect 1402 3143 1413 3146
rect 1410 3133 1413 3143
rect 1410 3033 1413 3126
rect 1418 3096 1421 3153
rect 1434 3133 1437 3176
rect 1442 3146 1445 3216
rect 1462 3146 1465 3223
rect 1442 3143 1453 3146
rect 1458 3143 1465 3146
rect 1474 3213 1493 3216
rect 1458 3116 1461 3143
rect 1450 3113 1461 3116
rect 1418 3093 1429 3096
rect 1338 3023 1365 3026
rect 1394 3023 1405 3026
rect 1426 3023 1429 3093
rect 1450 3066 1453 3113
rect 1466 3073 1469 3126
rect 1474 3123 1477 3213
rect 1490 3176 1493 3213
rect 1530 3183 1533 3206
rect 1578 3176 1581 3216
rect 1490 3173 1517 3176
rect 1578 3173 1613 3176
rect 1490 3133 1493 3146
rect 1498 3133 1501 3146
rect 1482 3123 1493 3126
rect 1514 3123 1517 3173
rect 1482 3106 1485 3123
rect 1478 3103 1485 3106
rect 1490 3103 1493 3116
rect 1450 3063 1461 3066
rect 1322 2993 1325 3006
rect 1330 2973 1333 3006
rect 1266 2943 1285 2946
rect 1162 2913 1165 2936
rect 1170 2906 1173 2936
rect 1178 2923 1181 2936
rect 1186 2933 1205 2936
rect 1186 2913 1189 2933
rect 1170 2903 1189 2906
rect 1194 2896 1197 2926
rect 1162 2893 1197 2896
rect 1202 2893 1205 2933
rect 1210 2933 1221 2936
rect 1162 2836 1165 2893
rect 1162 2833 1173 2836
rect 962 2773 973 2776
rect 914 2623 917 2636
rect 922 2613 925 2646
rect 906 2603 917 2606
rect 890 2583 901 2586
rect 890 2556 893 2583
rect 898 2573 909 2576
rect 890 2553 897 2556
rect 894 2466 897 2553
rect 906 2523 909 2573
rect 930 2563 933 2666
rect 938 2613 941 2636
rect 946 2603 949 2626
rect 954 2613 957 2726
rect 962 2713 965 2773
rect 978 2753 989 2756
rect 978 2736 981 2753
rect 970 2733 981 2736
rect 970 2623 973 2733
rect 978 2693 981 2726
rect 986 2703 989 2736
rect 994 2723 997 2746
rect 1002 2696 1005 2766
rect 1034 2733 1053 2736
rect 1058 2733 1061 2756
rect 1050 2726 1053 2733
rect 1066 2726 1069 2736
rect 1090 2733 1093 2746
rect 1042 2713 1045 2726
rect 1050 2723 1061 2726
rect 1066 2723 1093 2726
rect 986 2693 1005 2696
rect 930 2533 933 2546
rect 938 2533 941 2576
rect 914 2476 917 2526
rect 954 2513 957 2606
rect 986 2586 989 2693
rect 994 2623 1037 2626
rect 994 2613 997 2623
rect 982 2583 989 2586
rect 970 2523 973 2556
rect 982 2526 985 2583
rect 994 2533 997 2576
rect 1002 2546 1005 2616
rect 1010 2613 1021 2616
rect 1010 2563 1013 2606
rect 1026 2603 1029 2616
rect 1034 2613 1037 2623
rect 1026 2566 1029 2586
rect 1026 2563 1033 2566
rect 1002 2543 1021 2546
rect 982 2523 989 2526
rect 914 2473 957 2476
rect 894 2463 925 2466
rect 874 2453 885 2456
rect 826 2403 829 2416
rect 810 2323 813 2336
rect 842 2323 845 2406
rect 874 2386 877 2453
rect 874 2383 885 2386
rect 882 2366 885 2383
rect 890 2376 893 2416
rect 922 2413 925 2463
rect 946 2406 949 2466
rect 954 2413 957 2473
rect 986 2463 989 2523
rect 1010 2483 1013 2536
rect 1018 2523 1021 2543
rect 1030 2516 1033 2563
rect 1042 2533 1045 2656
rect 1058 2616 1061 2716
rect 1090 2616 1093 2716
rect 1098 2713 1101 2736
rect 1106 2723 1109 2806
rect 1098 2633 1117 2636
rect 1098 2623 1101 2633
rect 1050 2613 1061 2616
rect 1026 2513 1033 2516
rect 946 2403 957 2406
rect 930 2383 933 2396
rect 890 2373 949 2376
rect 882 2363 893 2366
rect 858 2323 861 2346
rect 890 2323 893 2363
rect 770 2213 773 2226
rect 786 2213 789 2266
rect 802 2216 805 2286
rect 802 2213 821 2216
rect 778 2203 789 2206
rect 762 2193 789 2196
rect 794 2193 797 2206
rect 738 2173 749 2176
rect 714 2163 725 2166
rect 722 2146 725 2163
rect 698 2123 701 2136
rect 714 2133 717 2146
rect 722 2143 729 2146
rect 714 2106 717 2126
rect 706 2103 717 2106
rect 706 2056 709 2103
rect 706 2053 717 2056
rect 674 2023 701 2026
rect 666 2016 669 2023
rect 642 1963 653 1966
rect 618 1933 625 1936
rect 594 1763 597 1896
rect 570 1753 597 1756
rect 602 1753 605 1806
rect 610 1763 613 1816
rect 594 1746 597 1753
rect 562 1743 581 1746
rect 538 1613 541 1686
rect 546 1603 549 1736
rect 555 1723 565 1726
rect 570 1723 573 1736
rect 578 1723 581 1743
rect 546 1533 549 1556
rect 538 1523 549 1526
rect 538 1433 541 1466
rect 522 1416 525 1426
rect 530 1423 541 1426
rect 514 1403 517 1416
rect 522 1413 533 1416
rect 522 1383 525 1406
rect 538 1396 541 1423
rect 530 1393 541 1396
rect 530 1376 533 1393
rect 514 1373 533 1376
rect 514 1333 517 1373
rect 498 1323 517 1326
rect 498 943 501 1316
rect 490 933 501 936
rect 490 903 493 916
rect 490 803 493 866
rect 498 843 501 916
rect 498 773 501 816
rect 506 756 509 1296
rect 514 1213 517 1316
rect 522 1293 525 1336
rect 530 1233 533 1366
rect 538 1346 541 1386
rect 546 1353 549 1426
rect 538 1343 549 1346
rect 538 1296 541 1336
rect 546 1313 549 1343
rect 538 1293 549 1296
rect 538 1223 541 1256
rect 522 1213 541 1216
rect 546 1206 549 1293
rect 514 1153 517 1206
rect 538 1203 549 1206
rect 554 1203 557 1716
rect 562 1703 565 1723
rect 570 1713 581 1716
rect 570 1676 573 1713
rect 570 1673 581 1676
rect 562 1623 565 1636
rect 562 1573 565 1616
rect 562 1433 565 1566
rect 562 1413 565 1426
rect 570 1406 573 1666
rect 578 1583 581 1673
rect 578 1523 581 1576
rect 578 1423 581 1446
rect 562 1303 565 1406
rect 570 1403 577 1406
rect 574 1336 577 1403
rect 570 1333 577 1336
rect 562 1216 565 1286
rect 570 1263 573 1333
rect 562 1213 573 1216
rect 514 1063 517 1136
rect 522 1056 525 1146
rect 530 1113 533 1166
rect 538 1063 541 1203
rect 546 1173 557 1176
rect 522 1053 541 1056
rect 514 1003 525 1006
rect 530 1003 533 1026
rect 522 913 525 956
rect 538 946 541 1053
rect 546 953 549 1136
rect 554 1123 557 1173
rect 562 1116 565 1176
rect 570 1123 573 1213
rect 578 1203 581 1316
rect 586 1283 589 1746
rect 594 1743 605 1746
rect 594 1713 597 1736
rect 594 1563 597 1686
rect 602 1663 605 1743
rect 602 1633 605 1656
rect 594 1373 597 1536
rect 602 1533 605 1546
rect 610 1523 613 1726
rect 602 1413 605 1516
rect 610 1433 613 1476
rect 618 1463 621 1933
rect 634 1916 637 1936
rect 626 1913 637 1916
rect 626 1873 629 1913
rect 626 1823 629 1846
rect 626 1683 629 1806
rect 634 1803 637 1906
rect 642 1736 645 1956
rect 650 1893 653 1963
rect 658 1953 661 2016
rect 666 2013 685 2016
rect 698 2013 701 2023
rect 666 1996 669 2006
rect 682 1996 685 2006
rect 666 1993 685 1996
rect 666 1946 669 1986
rect 690 1983 693 2006
rect 658 1943 669 1946
rect 666 1923 677 1926
rect 658 1913 669 1916
rect 634 1733 645 1736
rect 634 1713 637 1726
rect 626 1623 629 1666
rect 626 1543 629 1616
rect 626 1446 629 1536
rect 634 1473 637 1636
rect 642 1613 645 1716
rect 650 1713 653 1886
rect 650 1606 653 1656
rect 642 1603 653 1606
rect 642 1533 645 1586
rect 618 1443 629 1446
rect 618 1426 621 1443
rect 610 1423 621 1426
rect 602 1356 605 1406
rect 610 1403 613 1423
rect 642 1416 645 1496
rect 650 1423 653 1516
rect 610 1363 613 1396
rect 594 1353 605 1356
rect 594 1296 597 1353
rect 618 1346 621 1416
rect 626 1413 636 1416
rect 642 1413 653 1416
rect 626 1403 629 1413
rect 602 1343 621 1346
rect 602 1323 605 1343
rect 610 1303 613 1336
rect 626 1333 629 1376
rect 618 1313 621 1326
rect 594 1293 613 1296
rect 578 1123 581 1196
rect 586 1163 589 1236
rect 554 1113 565 1116
rect 530 933 533 946
rect 538 943 549 946
rect 546 933 549 943
rect 530 916 533 926
rect 530 913 541 916
rect 514 893 517 906
rect 514 803 517 816
rect 522 796 525 826
rect 482 753 509 756
rect 514 793 525 796
rect 482 636 485 753
rect 498 733 501 746
rect 506 726 509 736
rect 514 733 517 793
rect 530 776 533 896
rect 526 773 533 776
rect 490 663 493 726
rect 506 723 517 726
rect 474 633 485 636
rect 458 613 461 626
rect 474 606 477 633
rect 482 613 485 626
rect 498 623 501 676
rect 466 603 477 606
rect 442 583 449 586
rect 430 503 437 506
rect 430 436 433 503
rect 446 496 449 583
rect 466 546 469 603
rect 442 493 449 496
rect 458 543 469 546
rect 430 433 437 436
rect 394 383 405 386
rect 426 383 429 416
rect 434 396 437 433
rect 442 413 445 493
rect 442 403 453 406
rect 450 396 453 403
rect 458 396 461 543
rect 466 506 469 526
rect 490 513 493 536
rect 498 523 501 606
rect 466 503 477 506
rect 474 436 477 503
rect 434 393 445 396
rect 450 393 461 396
rect 470 433 477 436
rect 402 376 405 383
rect 402 373 437 376
rect 402 323 405 373
rect 374 313 381 316
rect 258 213 269 216
rect 258 203 261 213
rect 274 193 277 226
rect 282 213 285 226
rect 274 123 277 136
rect 282 123 285 166
rect 306 146 309 283
rect 322 236 325 303
rect 378 256 381 313
rect 402 313 421 316
rect 426 313 429 366
rect 434 323 437 373
rect 442 316 445 393
rect 470 386 473 433
rect 466 383 473 386
rect 466 326 469 383
rect 466 323 473 326
rect 434 313 445 316
rect 378 253 389 256
rect 318 233 325 236
rect 318 166 321 233
rect 362 226 365 236
rect 330 223 365 226
rect 318 163 325 166
rect 306 143 317 146
rect 314 123 317 143
rect 322 133 325 163
rect 330 123 333 223
rect 338 123 341 196
rect 346 186 349 206
rect 354 196 357 216
rect 362 203 365 223
rect 370 213 373 246
rect 370 196 373 206
rect 354 193 373 196
rect 386 186 389 253
rect 346 183 389 186
rect 346 143 373 146
rect 346 133 349 143
rect 354 123 357 136
rect 370 133 373 143
rect 90 103 97 106
rect 90 83 93 103
rect 362 93 365 126
rect 386 123 389 136
rect 402 133 405 313
rect 410 296 413 306
rect 426 296 429 306
rect 410 293 429 296
rect 410 213 421 216
rect 434 213 437 313
rect 442 146 445 226
rect 450 213 453 256
rect 458 233 461 316
rect 470 226 473 323
rect 482 263 485 416
rect 498 366 501 406
rect 490 363 501 366
rect 506 363 509 723
rect 514 586 517 696
rect 526 636 529 773
rect 526 633 533 636
rect 522 603 525 616
rect 530 593 533 633
rect 514 583 533 586
rect 514 533 525 536
rect 514 513 517 533
rect 530 493 533 583
rect 514 413 517 426
rect 538 406 541 913
rect 546 413 549 906
rect 554 843 557 1113
rect 554 813 557 826
rect 562 786 565 1106
rect 578 1066 581 1116
rect 586 1073 589 1136
rect 578 1063 589 1066
rect 570 993 573 1016
rect 570 923 573 966
rect 570 863 573 906
rect 578 813 581 1026
rect 586 983 589 1063
rect 594 1033 597 1226
rect 602 1213 605 1226
rect 602 1083 605 1206
rect 610 1203 613 1293
rect 618 1196 621 1236
rect 626 1223 629 1276
rect 610 1193 621 1196
rect 610 1016 613 1193
rect 618 1096 621 1146
rect 626 1103 629 1136
rect 618 1093 625 1096
rect 622 1036 625 1093
rect 622 1033 629 1036
rect 594 1003 597 1016
rect 602 1013 621 1016
rect 602 976 605 1013
rect 586 973 605 976
rect 586 903 589 973
rect 594 956 597 966
rect 610 963 613 1006
rect 618 1003 621 1013
rect 594 953 621 956
rect 610 926 613 936
rect 594 893 597 926
rect 602 923 613 926
rect 570 803 581 806
rect 554 783 565 786
rect 514 403 541 406
rect 554 396 557 783
rect 562 623 565 726
rect 570 686 573 736
rect 578 723 581 776
rect 586 703 589 836
rect 594 803 597 816
rect 602 796 605 923
rect 610 813 613 916
rect 618 806 621 936
rect 626 863 629 1033
rect 634 953 637 1366
rect 642 1306 645 1406
rect 650 1323 653 1413
rect 658 1323 661 1906
rect 666 1843 669 1913
rect 674 1893 677 1923
rect 682 1903 685 1956
rect 666 1806 669 1826
rect 674 1813 677 1876
rect 682 1813 685 1886
rect 666 1803 677 1806
rect 690 1796 693 1926
rect 698 1916 701 2006
rect 714 1983 717 2053
rect 726 2026 729 2143
rect 746 2116 749 2173
rect 738 2113 749 2116
rect 738 2093 741 2113
rect 722 2023 729 2026
rect 706 1943 709 1956
rect 714 1933 717 1946
rect 722 1923 725 2023
rect 730 1946 733 2006
rect 738 2003 741 2036
rect 762 2013 765 2066
rect 770 2016 773 2136
rect 786 2133 789 2193
rect 802 2143 805 2206
rect 778 2063 781 2126
rect 794 2076 797 2136
rect 810 2133 813 2206
rect 818 2196 821 2213
rect 818 2193 829 2196
rect 826 2146 829 2193
rect 842 2153 845 2226
rect 818 2143 829 2146
rect 818 2126 821 2143
rect 786 2073 797 2076
rect 802 2073 805 2126
rect 810 2123 821 2126
rect 770 2013 781 2016
rect 786 2013 789 2073
rect 754 1973 757 2006
rect 730 1943 757 1946
rect 738 1926 741 1936
rect 730 1923 741 1926
rect 698 1913 709 1916
rect 730 1913 733 1923
rect 674 1793 693 1796
rect 674 1733 677 1793
rect 666 1713 677 1716
rect 666 1623 669 1666
rect 682 1636 685 1666
rect 674 1633 685 1636
rect 666 1583 669 1606
rect 674 1526 677 1633
rect 682 1603 685 1626
rect 690 1613 693 1766
rect 698 1733 701 1846
rect 706 1836 709 1913
rect 738 1906 741 1916
rect 722 1903 741 1906
rect 706 1833 713 1836
rect 710 1756 713 1833
rect 706 1753 713 1756
rect 698 1713 701 1726
rect 706 1663 709 1753
rect 698 1623 709 1626
rect 698 1596 701 1623
rect 666 1523 677 1526
rect 666 1373 669 1523
rect 682 1486 685 1596
rect 698 1593 709 1596
rect 690 1533 693 1586
rect 674 1483 685 1486
rect 674 1443 677 1483
rect 690 1476 693 1506
rect 682 1473 693 1476
rect 682 1413 685 1473
rect 690 1403 693 1466
rect 698 1423 701 1576
rect 706 1523 709 1593
rect 698 1386 701 1416
rect 694 1383 701 1386
rect 666 1323 669 1336
rect 642 1303 649 1306
rect 646 1246 649 1303
rect 658 1253 661 1316
rect 646 1243 661 1246
rect 666 1243 669 1316
rect 674 1303 677 1366
rect 694 1316 697 1383
rect 682 1303 685 1316
rect 694 1313 701 1316
rect 674 1293 693 1296
rect 642 1133 645 1206
rect 650 1123 653 1216
rect 642 1013 645 1026
rect 642 993 645 1006
rect 650 1003 653 1056
rect 658 996 661 1243
rect 666 1123 669 1226
rect 666 1023 669 1086
rect 650 993 661 996
rect 626 813 629 836
rect 598 793 605 796
rect 610 793 613 806
rect 618 803 629 806
rect 598 736 601 793
rect 594 733 601 736
rect 610 733 613 746
rect 594 713 597 733
rect 570 683 597 686
rect 570 613 573 636
rect 562 593 565 606
rect 562 513 565 586
rect 586 553 589 616
rect 594 613 597 683
rect 618 633 621 756
rect 626 723 629 803
rect 634 633 637 906
rect 618 603 621 616
rect 586 523 597 526
rect 602 523 605 536
rect 626 533 629 546
rect 602 513 621 516
rect 538 393 557 396
rect 490 316 493 363
rect 490 313 501 316
rect 522 313 525 336
rect 530 333 533 356
rect 538 326 541 393
rect 562 383 565 486
rect 602 406 605 513
rect 626 506 629 526
rect 610 503 629 506
rect 642 483 645 906
rect 650 803 653 993
rect 658 813 661 936
rect 658 796 661 806
rect 650 793 661 796
rect 650 733 653 793
rect 658 726 661 786
rect 650 723 661 726
rect 650 653 653 723
rect 666 666 669 956
rect 674 733 677 1293
rect 698 1273 701 1313
rect 706 1303 709 1486
rect 682 1193 685 1206
rect 682 1133 685 1156
rect 682 1056 685 1126
rect 690 1123 693 1216
rect 698 1173 701 1256
rect 706 1213 709 1296
rect 714 1186 717 1736
rect 722 1286 725 1903
rect 746 1896 749 1936
rect 754 1903 757 1943
rect 730 1893 761 1896
rect 730 1733 733 1893
rect 738 1806 741 1876
rect 746 1813 749 1836
rect 758 1826 761 1893
rect 758 1823 765 1826
rect 770 1823 773 2006
rect 778 1986 781 2013
rect 786 1993 789 2006
rect 810 1996 813 2123
rect 818 2003 821 2016
rect 826 2013 829 2116
rect 834 2003 837 2096
rect 794 1993 813 1996
rect 778 1983 789 1986
rect 794 1976 797 1993
rect 778 1973 797 1976
rect 778 1893 781 1973
rect 802 1943 805 1986
rect 810 1933 813 1946
rect 842 1943 845 2066
rect 850 2033 853 2206
rect 858 2146 861 2316
rect 874 2213 877 2226
rect 866 2173 869 2206
rect 882 2203 885 2286
rect 898 2213 901 2336
rect 914 2326 917 2356
rect 946 2333 949 2373
rect 954 2366 957 2403
rect 962 2376 965 2406
rect 978 2403 981 2456
rect 1010 2426 1013 2476
rect 1010 2423 1017 2426
rect 1002 2376 1005 2416
rect 962 2373 1005 2376
rect 1014 2366 1017 2423
rect 1026 2383 1029 2513
rect 1050 2506 1053 2613
rect 1074 2546 1077 2616
rect 1090 2613 1101 2616
rect 1106 2613 1109 2626
rect 1114 2616 1117 2633
rect 1122 2623 1125 2806
rect 1130 2723 1133 2816
rect 1170 2813 1173 2833
rect 1178 2803 1181 2886
rect 1138 2733 1141 2756
rect 1186 2746 1189 2846
rect 1210 2833 1213 2933
rect 1218 2903 1221 2926
rect 1226 2913 1229 2936
rect 1250 2913 1253 2936
rect 1258 2903 1261 2926
rect 1266 2876 1269 2943
rect 1274 2903 1277 2926
rect 1282 2893 1285 2926
rect 1290 2896 1293 2953
rect 1298 2906 1301 2936
rect 1338 2933 1341 3023
rect 1346 2976 1349 3006
rect 1354 2993 1357 3016
rect 1362 3013 1365 3023
rect 1370 3003 1373 3016
rect 1378 3013 1397 3016
rect 1394 2993 1397 3006
rect 1402 2983 1405 3023
rect 1410 2976 1413 3016
rect 1418 3013 1429 3016
rect 1458 3006 1461 3063
rect 1434 2983 1437 3006
rect 1442 2976 1445 3006
rect 1346 2973 1353 2976
rect 1410 2973 1445 2976
rect 1350 2926 1353 2973
rect 1442 2956 1445 2973
rect 1450 3003 1461 3006
rect 1450 2963 1453 3003
rect 1458 2973 1461 2996
rect 1442 2953 1453 2956
rect 1370 2943 1421 2946
rect 1306 2923 1317 2926
rect 1306 2913 1317 2916
rect 1322 2906 1325 2926
rect 1346 2923 1353 2926
rect 1298 2903 1317 2906
rect 1322 2903 1333 2906
rect 1290 2893 1325 2896
rect 1258 2873 1269 2876
rect 1250 2823 1253 2846
rect 1178 2743 1197 2746
rect 1138 2716 1141 2726
rect 1146 2723 1149 2736
rect 1138 2713 1157 2716
rect 1162 2713 1165 2736
rect 1178 2726 1181 2743
rect 1170 2723 1181 2726
rect 1170 2713 1189 2716
rect 1154 2703 1157 2713
rect 1170 2703 1173 2713
rect 1202 2706 1205 2796
rect 1178 2703 1205 2706
rect 1138 2623 1149 2626
rect 1162 2623 1165 2646
rect 1114 2613 1133 2616
rect 1146 2613 1149 2623
rect 1058 2533 1061 2546
rect 1074 2543 1085 2546
rect 1066 2523 1069 2536
rect 1050 2503 1061 2506
rect 1074 2483 1077 2536
rect 1082 2533 1085 2543
rect 1082 2503 1085 2526
rect 1090 2473 1093 2596
rect 1098 2533 1101 2613
rect 1130 2593 1133 2606
rect 1106 2533 1109 2556
rect 1114 2523 1117 2536
rect 1122 2533 1125 2576
rect 1074 2413 1077 2426
rect 954 2363 965 2366
rect 914 2323 925 2326
rect 922 2213 925 2323
rect 930 2203 933 2226
rect 858 2143 869 2146
rect 874 2143 885 2146
rect 858 2026 861 2136
rect 866 2063 869 2143
rect 874 2033 877 2136
rect 826 1933 845 1936
rect 802 1866 805 1926
rect 810 1913 813 1926
rect 778 1863 805 1866
rect 738 1803 757 1806
rect 738 1726 741 1736
rect 734 1723 741 1726
rect 734 1626 737 1723
rect 730 1623 737 1626
rect 730 1483 733 1623
rect 746 1613 749 1726
rect 754 1713 757 1803
rect 762 1703 765 1823
rect 770 1786 773 1816
rect 778 1803 781 1863
rect 810 1853 829 1856
rect 810 1826 813 1853
rect 786 1823 813 1826
rect 826 1823 829 1853
rect 850 1836 853 2026
rect 858 2023 877 2026
rect 858 1923 861 2006
rect 866 1983 869 1996
rect 866 1893 869 1946
rect 850 1833 861 1836
rect 818 1786 821 1806
rect 826 1803 829 1816
rect 770 1783 781 1786
rect 778 1696 781 1783
rect 810 1783 821 1786
rect 810 1736 813 1783
rect 810 1733 817 1736
rect 770 1693 781 1696
rect 770 1616 773 1693
rect 794 1626 797 1646
rect 790 1623 797 1626
rect 754 1613 781 1616
rect 738 1586 741 1606
rect 754 1603 757 1613
rect 738 1583 745 1586
rect 742 1516 745 1583
rect 738 1513 745 1516
rect 730 1413 733 1446
rect 730 1303 733 1406
rect 738 1363 741 1513
rect 746 1443 749 1496
rect 746 1346 749 1436
rect 738 1343 749 1346
rect 722 1283 729 1286
rect 706 1183 717 1186
rect 682 1053 693 1056
rect 682 903 685 1053
rect 698 1033 701 1136
rect 706 1066 709 1183
rect 714 1123 717 1176
rect 726 1166 729 1283
rect 738 1203 741 1343
rect 746 1233 749 1336
rect 746 1213 749 1226
rect 726 1163 733 1166
rect 722 1083 725 1126
rect 730 1076 733 1163
rect 738 1133 741 1156
rect 754 1143 757 1526
rect 762 1503 765 1566
rect 778 1536 781 1606
rect 790 1546 793 1623
rect 790 1543 797 1546
rect 770 1533 781 1536
rect 762 1173 765 1486
rect 770 1436 773 1466
rect 778 1446 781 1526
rect 794 1493 797 1543
rect 802 1533 805 1716
rect 814 1646 817 1733
rect 814 1643 821 1646
rect 778 1443 805 1446
rect 770 1433 789 1436
rect 770 1413 781 1416
rect 746 1133 757 1136
rect 738 1103 741 1126
rect 722 1073 733 1076
rect 706 1063 717 1066
rect 690 1003 701 1006
rect 706 996 709 1026
rect 698 993 709 996
rect 714 986 717 1063
rect 722 1016 725 1073
rect 730 1033 733 1056
rect 722 1013 729 1016
rect 682 796 685 836
rect 690 803 693 926
rect 698 913 701 986
rect 706 983 717 986
rect 698 863 701 906
rect 682 793 693 796
rect 682 733 685 776
rect 674 716 677 726
rect 690 723 693 793
rect 698 716 701 846
rect 706 766 709 983
rect 714 933 717 956
rect 726 936 729 1013
rect 722 933 729 936
rect 722 913 725 933
rect 738 906 741 1066
rect 746 1053 749 1126
rect 746 923 749 1036
rect 754 916 757 1133
rect 762 956 765 1136
rect 770 966 773 1406
rect 786 1373 789 1433
rect 794 1423 797 1436
rect 778 1223 781 1336
rect 786 1276 789 1356
rect 794 1313 797 1416
rect 802 1403 805 1443
rect 810 1336 813 1626
rect 818 1586 821 1643
rect 826 1603 829 1796
rect 850 1726 853 1826
rect 858 1736 861 1833
rect 866 1803 869 1816
rect 874 1773 877 2023
rect 882 1923 885 2066
rect 890 2003 893 2196
rect 898 2106 901 2166
rect 946 2163 949 2316
rect 954 2303 957 2336
rect 962 2256 965 2363
rect 1010 2363 1017 2366
rect 978 2333 981 2346
rect 978 2266 981 2316
rect 978 2263 985 2266
rect 962 2253 973 2256
rect 954 2146 957 2206
rect 962 2203 965 2236
rect 970 2213 973 2253
rect 982 2206 985 2263
rect 1010 2256 1013 2363
rect 1082 2336 1085 2416
rect 1090 2383 1093 2406
rect 1098 2366 1101 2486
rect 1114 2413 1117 2496
rect 1130 2483 1133 2546
rect 1138 2506 1141 2536
rect 1146 2513 1149 2606
rect 1178 2576 1181 2636
rect 1194 2576 1197 2676
rect 1210 2623 1213 2726
rect 1218 2723 1221 2816
rect 1258 2813 1261 2873
rect 1298 2803 1301 2816
rect 1322 2813 1325 2893
rect 1330 2873 1333 2903
rect 1346 2856 1349 2923
rect 1362 2903 1365 2916
rect 1342 2853 1349 2856
rect 1342 2796 1345 2853
rect 1226 2726 1229 2756
rect 1234 2733 1237 2746
rect 1226 2723 1237 2726
rect 1234 2706 1237 2723
rect 1226 2703 1237 2706
rect 1226 2636 1229 2703
rect 1226 2633 1237 2636
rect 1234 2613 1237 2633
rect 1242 2596 1245 2776
rect 1290 2743 1301 2746
rect 1250 2696 1253 2716
rect 1266 2713 1269 2736
rect 1322 2733 1325 2786
rect 1282 2723 1293 2726
rect 1250 2693 1261 2696
rect 1258 2636 1261 2693
rect 1170 2573 1181 2576
rect 1186 2573 1197 2576
rect 1170 2533 1173 2573
rect 1170 2506 1173 2526
rect 1138 2503 1173 2506
rect 1122 2413 1125 2436
rect 1138 2413 1141 2503
rect 1170 2473 1173 2503
rect 1178 2466 1181 2536
rect 1186 2523 1189 2573
rect 1202 2566 1205 2576
rect 1194 2563 1205 2566
rect 1218 2563 1221 2596
rect 1238 2593 1245 2596
rect 1250 2633 1261 2636
rect 1194 2533 1197 2563
rect 1194 2503 1197 2526
rect 1210 2513 1213 2536
rect 1218 2523 1221 2536
rect 1226 2506 1229 2536
rect 1202 2503 1229 2506
rect 1202 2466 1205 2503
rect 1238 2496 1241 2593
rect 1250 2503 1253 2633
rect 1258 2573 1261 2606
rect 1266 2593 1269 2606
rect 1282 2593 1285 2606
rect 1178 2463 1205 2466
rect 1162 2413 1165 2446
rect 1098 2363 1109 2366
rect 1042 2323 1045 2336
rect 1082 2333 1093 2336
rect 1090 2306 1093 2326
rect 1082 2303 1093 2306
rect 1010 2253 1021 2256
rect 978 2203 985 2206
rect 906 2143 917 2146
rect 930 2143 957 2146
rect 906 2113 909 2143
rect 898 2103 917 2106
rect 898 2043 901 2066
rect 890 1916 893 1986
rect 906 1973 909 2096
rect 914 2076 917 2103
rect 922 2083 925 2136
rect 914 2073 925 2076
rect 914 2013 917 2026
rect 914 1956 917 1986
rect 882 1913 893 1916
rect 898 1953 917 1956
rect 858 1733 869 1736
rect 842 1713 845 1726
rect 850 1723 861 1726
rect 850 1696 853 1716
rect 842 1693 853 1696
rect 842 1646 845 1693
rect 842 1643 853 1646
rect 850 1623 853 1643
rect 818 1583 825 1586
rect 822 1506 825 1583
rect 802 1333 813 1336
rect 818 1503 825 1506
rect 786 1273 797 1276
rect 778 1113 781 1216
rect 786 1203 789 1216
rect 794 1213 797 1273
rect 802 1206 805 1333
rect 810 1273 813 1326
rect 810 1213 813 1236
rect 794 1203 805 1206
rect 794 1133 797 1203
rect 802 1133 805 1196
rect 810 1133 813 1176
rect 794 1123 805 1126
rect 778 1013 781 1086
rect 778 993 781 1006
rect 770 963 781 966
rect 762 953 773 956
rect 770 933 773 953
rect 722 903 741 906
rect 746 913 757 916
rect 714 813 717 846
rect 722 833 725 903
rect 722 813 733 816
rect 722 783 725 806
rect 706 763 717 766
rect 674 713 701 716
rect 698 696 701 713
rect 658 663 669 666
rect 690 693 701 696
rect 650 623 653 636
rect 650 523 653 536
rect 618 423 645 426
rect 586 326 589 406
rect 602 403 613 406
rect 530 323 541 326
rect 498 256 501 313
rect 466 223 473 226
rect 490 253 501 256
rect 466 203 469 223
rect 442 143 453 146
rect 450 123 453 143
rect 466 123 469 146
rect 490 133 493 253
rect 522 223 525 236
rect 530 206 533 323
rect 546 213 549 326
rect 554 323 589 326
rect 594 316 597 396
rect 594 313 605 316
rect 610 296 613 403
rect 626 393 629 416
rect 642 413 645 423
rect 658 413 661 663
rect 666 503 669 656
rect 674 406 677 626
rect 690 616 693 693
rect 714 686 717 763
rect 706 683 717 686
rect 690 613 697 616
rect 682 543 685 596
rect 694 556 697 613
rect 706 593 709 683
rect 714 586 717 626
rect 730 613 733 736
rect 738 686 741 836
rect 746 696 749 913
rect 754 796 757 846
rect 762 803 765 926
rect 778 916 781 963
rect 774 913 781 916
rect 774 846 777 913
rect 774 843 781 846
rect 778 823 781 843
rect 754 793 765 796
rect 754 733 757 756
rect 754 706 757 726
rect 762 723 765 793
rect 770 733 773 746
rect 754 703 765 706
rect 746 693 769 696
rect 738 683 745 686
rect 706 583 717 586
rect 694 553 701 556
rect 690 516 693 536
rect 698 533 701 553
rect 686 513 693 516
rect 686 426 689 513
rect 698 433 701 526
rect 706 503 709 583
rect 686 423 693 426
rect 706 423 709 436
rect 634 386 637 406
rect 626 383 637 386
rect 642 403 653 406
rect 666 403 677 406
rect 602 293 613 296
rect 602 226 605 293
rect 618 243 621 336
rect 626 333 629 383
rect 642 336 645 403
rect 650 393 661 396
rect 658 376 661 393
rect 634 333 645 336
rect 654 373 661 376
rect 634 303 637 326
rect 654 316 657 373
rect 666 323 669 403
rect 674 333 677 386
rect 690 376 693 423
rect 714 413 717 536
rect 722 513 725 576
rect 730 436 733 606
rect 742 556 745 683
rect 742 553 749 556
rect 738 523 741 536
rect 746 496 749 553
rect 754 543 757 676
rect 766 626 769 693
rect 766 623 773 626
rect 762 593 765 606
rect 770 523 773 623
rect 778 613 781 816
rect 722 433 733 436
rect 742 493 749 496
rect 742 436 745 493
rect 742 433 749 436
rect 686 373 693 376
rect 674 316 677 326
rect 686 316 689 373
rect 698 323 701 366
rect 654 313 661 316
rect 674 313 689 316
rect 522 203 533 206
rect 522 146 525 203
rect 554 183 557 226
rect 602 223 613 226
rect 538 173 557 176
rect 522 143 533 146
rect 530 123 533 143
rect 538 133 541 173
rect 586 123 589 136
rect 594 123 597 206
rect 602 193 605 206
rect 610 133 613 223
rect 618 173 621 216
rect 626 213 637 216
rect 642 193 645 216
rect 658 203 661 313
rect 698 303 701 316
rect 706 286 709 336
rect 698 283 709 286
rect 682 246 685 266
rect 682 243 689 246
rect 674 203 677 226
rect 686 196 689 243
rect 698 236 701 283
rect 698 233 709 236
rect 706 213 709 233
rect 714 203 717 326
rect 722 223 725 433
rect 730 393 733 426
rect 738 326 741 416
rect 730 323 741 326
rect 682 193 689 196
rect 594 113 605 116
rect 602 76 605 113
rect 618 76 621 126
rect 634 123 637 146
rect 674 133 677 146
rect 682 133 685 193
rect 730 143 733 323
rect 738 223 741 316
rect 746 293 749 433
rect 754 403 757 486
rect 770 423 773 446
rect 770 333 773 406
rect 778 346 781 606
rect 786 433 789 1116
rect 794 1013 797 1116
rect 802 1073 805 1123
rect 810 1103 813 1126
rect 802 1006 805 1056
rect 818 1043 821 1503
rect 826 1126 829 1486
rect 834 1393 837 1596
rect 842 1433 845 1576
rect 850 1483 853 1606
rect 858 1603 861 1723
rect 866 1686 869 1733
rect 874 1703 877 1736
rect 866 1683 873 1686
rect 870 1596 873 1683
rect 866 1593 873 1596
rect 858 1533 861 1546
rect 834 1223 837 1386
rect 834 1133 837 1216
rect 842 1193 845 1426
rect 850 1343 853 1446
rect 850 1293 853 1336
rect 850 1213 853 1286
rect 858 1256 861 1406
rect 866 1393 869 1593
rect 874 1493 877 1526
rect 882 1406 885 1913
rect 898 1803 901 1953
rect 906 1923 909 1936
rect 914 1813 917 1886
rect 890 1733 893 1746
rect 898 1716 901 1796
rect 894 1713 901 1716
rect 894 1636 897 1713
rect 894 1633 901 1636
rect 890 1533 893 1556
rect 898 1536 901 1633
rect 906 1623 909 1746
rect 914 1713 917 1806
rect 906 1546 909 1616
rect 914 1583 917 1666
rect 906 1543 917 1546
rect 898 1533 909 1536
rect 890 1503 893 1526
rect 898 1493 901 1526
rect 878 1403 885 1406
rect 898 1406 901 1436
rect 906 1413 909 1533
rect 914 1483 917 1543
rect 914 1423 917 1456
rect 898 1403 909 1406
rect 922 1403 925 2073
rect 930 1823 933 2143
rect 938 2083 941 2136
rect 946 2133 957 2136
rect 946 2123 957 2126
rect 938 1913 941 2016
rect 946 2013 949 2116
rect 954 2093 957 2123
rect 946 1983 949 2006
rect 946 1943 949 1976
rect 938 1813 941 1896
rect 946 1806 949 1936
rect 954 1916 957 2046
rect 962 1993 965 2126
rect 962 1933 965 1966
rect 970 1933 973 2136
rect 954 1913 961 1916
rect 930 1743 933 1806
rect 938 1803 949 1806
rect 938 1646 941 1803
rect 958 1796 961 1913
rect 954 1793 961 1796
rect 954 1736 957 1793
rect 954 1733 965 1736
rect 954 1713 957 1726
rect 962 1663 965 1733
rect 930 1643 941 1646
rect 930 1433 933 1643
rect 938 1603 941 1626
rect 954 1613 965 1616
rect 878 1356 881 1403
rect 878 1353 885 1356
rect 866 1316 869 1336
rect 874 1323 877 1336
rect 882 1316 885 1353
rect 866 1313 885 1316
rect 858 1253 877 1256
rect 866 1226 869 1246
rect 862 1223 869 1226
rect 842 1133 845 1176
rect 826 1123 845 1126
rect 834 1086 837 1116
rect 826 1083 837 1086
rect 794 1003 805 1006
rect 810 1033 821 1036
rect 826 1033 829 1083
rect 842 1076 845 1123
rect 834 1073 845 1076
rect 794 806 797 1003
rect 802 943 805 956
rect 810 933 813 1033
rect 818 983 821 1026
rect 818 933 821 956
rect 802 813 805 916
rect 818 906 821 926
rect 814 903 821 906
rect 814 836 817 903
rect 814 833 821 836
rect 818 813 821 833
rect 794 803 805 806
rect 794 703 797 736
rect 802 696 805 803
rect 794 693 805 696
rect 810 803 821 806
rect 786 403 789 426
rect 778 343 785 346
rect 754 323 773 326
rect 754 303 757 323
rect 762 236 765 316
rect 770 313 773 323
rect 782 286 785 343
rect 782 283 789 286
rect 786 266 789 283
rect 778 263 789 266
rect 754 233 765 236
rect 794 233 797 693
rect 802 393 805 686
rect 810 613 813 803
rect 818 643 821 726
rect 826 613 829 1026
rect 834 993 837 1073
rect 842 1013 845 1066
rect 834 796 837 986
rect 842 936 845 1006
rect 850 1003 853 1206
rect 862 1146 865 1223
rect 862 1143 869 1146
rect 858 1016 861 1126
rect 866 1033 869 1143
rect 874 1053 877 1253
rect 882 1203 885 1313
rect 890 1303 893 1396
rect 882 1093 885 1196
rect 890 1166 893 1216
rect 898 1173 901 1336
rect 906 1166 909 1403
rect 930 1336 933 1426
rect 938 1403 941 1586
rect 946 1396 949 1486
rect 954 1413 957 1556
rect 962 1473 965 1606
rect 962 1423 965 1456
rect 914 1303 917 1336
rect 922 1333 933 1336
rect 938 1393 949 1396
rect 890 1163 909 1166
rect 914 1146 917 1206
rect 922 1193 925 1333
rect 938 1326 941 1393
rect 934 1323 941 1326
rect 934 1246 937 1323
rect 930 1243 937 1246
rect 930 1186 933 1243
rect 946 1226 949 1366
rect 938 1223 949 1226
rect 910 1143 917 1146
rect 922 1183 933 1186
rect 858 1013 869 1016
rect 850 946 853 996
rect 858 953 861 1006
rect 866 956 869 1013
rect 874 993 877 1016
rect 882 1003 885 1066
rect 890 1036 893 1086
rect 898 1043 901 1136
rect 910 1086 913 1143
rect 922 1093 925 1183
rect 938 1133 941 1206
rect 946 1133 949 1216
rect 910 1083 917 1086
rect 914 1066 917 1083
rect 906 1063 917 1066
rect 890 1033 909 1036
rect 890 1013 893 1026
rect 898 986 901 1026
rect 906 1003 909 1033
rect 890 983 901 986
rect 866 953 877 956
rect 850 943 869 946
rect 842 933 853 936
rect 842 913 845 926
rect 842 803 845 826
rect 834 793 845 796
rect 850 793 853 896
rect 858 803 861 936
rect 866 893 869 943
rect 874 893 877 953
rect 890 886 893 983
rect 890 883 901 886
rect 810 593 813 606
rect 834 596 837 786
rect 842 683 845 793
rect 818 593 837 596
rect 810 523 813 536
rect 818 496 821 593
rect 842 573 845 606
rect 850 603 853 736
rect 858 733 861 796
rect 858 703 861 716
rect 826 533 837 536
rect 826 513 829 526
rect 842 523 845 536
rect 850 533 853 556
rect 858 533 861 616
rect 850 523 861 526
rect 810 326 813 496
rect 818 493 829 496
rect 826 426 829 493
rect 818 423 829 426
rect 818 403 821 423
rect 842 376 845 416
rect 850 403 853 436
rect 858 423 861 446
rect 834 373 845 376
rect 802 323 813 326
rect 754 216 757 233
rect 750 213 757 216
rect 762 223 813 226
rect 818 223 821 336
rect 834 326 837 373
rect 850 333 853 366
rect 834 323 845 326
rect 750 156 753 213
rect 750 153 757 156
rect 690 133 701 136
rect 698 113 701 126
rect 738 123 741 136
rect 754 133 757 153
rect 746 103 749 126
rect 762 123 765 223
rect 786 166 789 206
rect 794 193 797 206
rect 786 163 797 166
rect 602 73 621 76
rect 778 53 781 156
rect 794 96 797 163
rect 810 133 813 216
rect 842 203 845 323
rect 858 313 861 416
rect 866 296 869 816
rect 874 723 877 836
rect 882 636 885 866
rect 874 633 885 636
rect 874 583 877 626
rect 874 433 877 536
rect 882 533 885 616
rect 890 423 893 846
rect 898 793 901 883
rect 898 703 901 726
rect 906 706 909 986
rect 914 723 917 1056
rect 922 796 925 1036
rect 930 983 933 1126
rect 930 923 933 946
rect 930 813 933 846
rect 922 793 929 796
rect 926 716 929 793
rect 922 713 929 716
rect 906 703 913 706
rect 898 586 901 676
rect 910 606 913 703
rect 922 623 925 713
rect 910 603 917 606
rect 930 603 933 646
rect 898 583 905 586
rect 902 496 905 583
rect 898 493 905 496
rect 898 473 901 493
rect 914 466 917 603
rect 930 523 933 536
rect 938 516 941 1086
rect 946 1063 949 1126
rect 946 993 949 1016
rect 946 893 949 936
rect 946 783 949 816
rect 946 693 949 736
rect 954 673 957 1406
rect 962 1373 965 1396
rect 962 1203 965 1336
rect 970 1246 973 1866
rect 978 1453 981 2203
rect 994 2146 997 2226
rect 1002 2193 1005 2246
rect 1018 2166 1021 2253
rect 1034 2183 1037 2206
rect 1010 2163 1021 2166
rect 994 2143 1005 2146
rect 994 2123 997 2136
rect 986 2053 989 2116
rect 994 2013 997 2116
rect 1002 2043 1005 2143
rect 1010 2056 1013 2163
rect 1018 2073 1021 2126
rect 1010 2053 1017 2056
rect 986 1933 989 1956
rect 994 1923 997 1996
rect 1002 1993 1005 2006
rect 1014 1976 1017 2053
rect 1026 2043 1029 2146
rect 1042 2133 1045 2296
rect 1082 2236 1085 2303
rect 1050 2086 1053 2226
rect 1058 2106 1061 2236
rect 1082 2233 1093 2236
rect 1074 2206 1077 2216
rect 1074 2203 1085 2206
rect 1090 2183 1093 2233
rect 1098 2203 1101 2256
rect 1106 2213 1109 2363
rect 1114 2306 1117 2396
rect 1122 2376 1125 2406
rect 1130 2383 1133 2406
rect 1146 2376 1149 2406
rect 1122 2373 1149 2376
rect 1146 2353 1149 2373
rect 1154 2363 1157 2406
rect 1122 2323 1125 2336
rect 1154 2323 1157 2336
rect 1114 2303 1125 2306
rect 1122 2236 1125 2303
rect 1114 2233 1125 2236
rect 1082 2123 1085 2166
rect 1106 2143 1109 2196
rect 1066 2113 1085 2116
rect 1082 2106 1085 2113
rect 1098 2106 1101 2116
rect 1106 2113 1109 2136
rect 1058 2103 1077 2106
rect 1082 2103 1101 2106
rect 1026 2003 1029 2026
rect 1034 2013 1037 2056
rect 1010 1973 1017 1976
rect 986 1723 989 1826
rect 994 1813 997 1916
rect 994 1703 997 1806
rect 986 1613 989 1646
rect 994 1613 997 1626
rect 986 1483 989 1606
rect 994 1533 997 1586
rect 1002 1553 1005 1956
rect 1010 1913 1013 1973
rect 1018 1906 1021 1956
rect 1014 1903 1021 1906
rect 1014 1826 1017 1903
rect 1010 1823 1017 1826
rect 1010 1803 1013 1823
rect 1026 1803 1029 1926
rect 1034 1916 1037 2006
rect 1042 1953 1045 2086
rect 1050 2083 1061 2086
rect 1058 1976 1061 2083
rect 1050 1973 1061 1976
rect 1050 1953 1053 1973
rect 1042 1943 1069 1946
rect 1042 1933 1045 1943
rect 1050 1933 1061 1936
rect 1066 1933 1069 1943
rect 1034 1913 1041 1916
rect 1038 1816 1041 1913
rect 1038 1813 1045 1816
rect 1002 1533 1005 1546
rect 1010 1533 1013 1766
rect 1034 1746 1037 1806
rect 1018 1743 1037 1746
rect 994 1483 997 1526
rect 978 1383 981 1426
rect 994 1376 997 1386
rect 978 1373 997 1376
rect 978 1343 981 1373
rect 1002 1356 1005 1466
rect 1010 1403 1013 1526
rect 1018 1443 1021 1743
rect 1042 1736 1045 1813
rect 1050 1803 1053 1926
rect 1058 1903 1061 1933
rect 1074 1836 1077 2103
rect 1082 2003 1085 2026
rect 1090 1883 1093 2066
rect 1098 1983 1101 2016
rect 1098 1903 1101 1926
rect 1106 1873 1109 2106
rect 1114 1986 1117 2233
rect 1122 2176 1125 2216
rect 1146 2213 1157 2216
rect 1130 2203 1141 2206
rect 1130 2183 1133 2203
rect 1122 2173 1137 2176
rect 1134 2126 1137 2173
rect 1146 2133 1149 2206
rect 1122 2103 1125 2126
rect 1134 2123 1141 2126
rect 1122 2003 1125 2036
rect 1130 2006 1133 2056
rect 1138 2013 1141 2123
rect 1154 2036 1157 2213
rect 1162 2183 1165 2246
rect 1170 2176 1173 2226
rect 1178 2206 1181 2346
rect 1186 2333 1189 2416
rect 1194 2326 1197 2416
rect 1202 2383 1205 2463
rect 1210 2366 1213 2446
rect 1218 2403 1221 2416
rect 1226 2413 1229 2496
rect 1238 2493 1245 2496
rect 1242 2443 1245 2493
rect 1266 2483 1269 2536
rect 1290 2533 1293 2723
rect 1314 2713 1317 2726
rect 1330 2676 1333 2796
rect 1342 2793 1349 2796
rect 1346 2776 1349 2793
rect 1346 2773 1357 2776
rect 1338 2723 1349 2726
rect 1322 2673 1333 2676
rect 1306 2613 1309 2646
rect 1298 2586 1301 2606
rect 1298 2583 1305 2586
rect 1302 2526 1305 2583
rect 1322 2576 1325 2673
rect 1354 2666 1357 2773
rect 1362 2733 1365 2776
rect 1338 2663 1357 2666
rect 1322 2573 1333 2576
rect 1298 2523 1305 2526
rect 1298 2476 1301 2523
rect 1314 2503 1317 2526
rect 1330 2486 1333 2573
rect 1338 2556 1341 2663
rect 1370 2656 1373 2866
rect 1378 2843 1381 2936
rect 1386 2883 1389 2926
rect 1394 2913 1397 2936
rect 1418 2933 1421 2943
rect 1402 2873 1405 2926
rect 1426 2923 1429 2946
rect 1434 2943 1445 2946
rect 1434 2933 1437 2943
rect 1450 2936 1453 2953
rect 1442 2933 1453 2936
rect 1442 2923 1445 2933
rect 1458 2926 1461 2936
rect 1450 2923 1461 2926
rect 1450 2916 1453 2923
rect 1426 2913 1453 2916
rect 1466 2913 1469 3016
rect 1478 2946 1481 3103
rect 1490 3003 1493 3096
rect 1522 3093 1525 3136
rect 1546 3106 1549 3126
rect 1554 3113 1565 3116
rect 1546 3103 1565 3106
rect 1570 3103 1573 3136
rect 1586 3133 1589 3166
rect 1610 3133 1613 3173
rect 1618 3133 1621 3146
rect 1634 3126 1637 3216
rect 1658 3183 1661 3206
rect 1706 3176 1709 3216
rect 1706 3173 1725 3176
rect 1594 3123 1637 3126
rect 1658 3116 1661 3136
rect 1682 3133 1685 3146
rect 1698 3133 1701 3166
rect 1722 3133 1725 3173
rect 1730 3133 1733 3146
rect 1738 3143 1741 3216
rect 1762 3183 1765 3206
rect 1794 3196 1797 3243
rect 1786 3193 1797 3196
rect 1786 3136 1789 3193
rect 1706 3123 1749 3126
rect 1474 2943 1481 2946
rect 1474 2906 1477 2943
rect 1498 2926 1501 3056
rect 1522 3023 1549 3026
rect 1522 3013 1525 3023
rect 1506 2993 1509 3006
rect 1522 2983 1525 3006
rect 1538 2996 1541 3016
rect 1546 3006 1549 3023
rect 1554 3013 1557 3036
rect 1546 3003 1557 3006
rect 1562 3003 1565 3103
rect 1570 3013 1573 3056
rect 1578 2996 1581 3006
rect 1538 2993 1581 2996
rect 1578 2983 1581 2993
rect 1482 2913 1485 2926
rect 1490 2916 1493 2926
rect 1498 2923 1509 2926
rect 1490 2913 1501 2916
rect 1466 2893 1469 2906
rect 1474 2903 1493 2906
rect 1378 2723 1381 2816
rect 1386 2713 1389 2806
rect 1402 2766 1405 2816
rect 1418 2793 1421 2816
rect 1450 2813 1453 2826
rect 1426 2773 1429 2806
rect 1466 2803 1469 2816
rect 1490 2813 1493 2903
rect 1498 2873 1501 2913
rect 1506 2793 1509 2923
rect 1514 2913 1517 2956
rect 1522 2903 1525 2926
rect 1538 2923 1541 2976
rect 1586 2973 1589 2996
rect 1554 2846 1557 2966
rect 1554 2843 1561 2846
rect 1546 2813 1549 2826
rect 1402 2763 1445 2766
rect 1442 2746 1445 2763
rect 1442 2743 1449 2746
rect 1346 2653 1373 2656
rect 1346 2576 1349 2653
rect 1362 2603 1365 2616
rect 1346 2573 1357 2576
rect 1338 2553 1345 2556
rect 1342 2486 1345 2553
rect 1202 2363 1213 2366
rect 1202 2353 1205 2363
rect 1186 2323 1197 2326
rect 1186 2303 1189 2323
rect 1202 2303 1205 2326
rect 1234 2323 1237 2436
rect 1242 2323 1245 2406
rect 1258 2363 1261 2406
rect 1274 2403 1277 2416
rect 1194 2213 1197 2286
rect 1202 2216 1205 2236
rect 1218 2216 1221 2276
rect 1258 2266 1261 2356
rect 1226 2263 1261 2266
rect 1226 2253 1229 2263
rect 1242 2233 1245 2256
rect 1258 2226 1261 2246
rect 1234 2223 1261 2226
rect 1202 2213 1209 2216
rect 1218 2213 1237 2216
rect 1178 2203 1197 2206
rect 1162 2173 1173 2176
rect 1162 2133 1165 2173
rect 1170 2093 1173 2126
rect 1154 2033 1173 2036
rect 1162 2016 1165 2026
rect 1154 2013 1165 2016
rect 1130 2003 1141 2006
rect 1114 1983 1125 1986
rect 1122 1866 1125 1983
rect 1138 1923 1141 2003
rect 1154 1953 1157 2013
rect 1138 1893 1141 1916
rect 1114 1863 1125 1866
rect 1066 1833 1085 1836
rect 1026 1733 1045 1736
rect 1026 1486 1029 1733
rect 1050 1726 1053 1776
rect 1034 1723 1053 1726
rect 1034 1656 1037 1716
rect 1034 1653 1045 1656
rect 1034 1523 1037 1646
rect 1042 1566 1045 1653
rect 1050 1633 1053 1723
rect 1058 1623 1061 1716
rect 1050 1603 1053 1616
rect 1066 1606 1069 1833
rect 1074 1796 1077 1826
rect 1082 1813 1085 1833
rect 1074 1793 1085 1796
rect 1082 1716 1085 1793
rect 1106 1786 1109 1806
rect 1078 1713 1085 1716
rect 1098 1783 1109 1786
rect 1078 1606 1081 1713
rect 1090 1613 1093 1646
rect 1062 1603 1069 1606
rect 1074 1603 1081 1606
rect 1050 1583 1053 1596
rect 1042 1563 1053 1566
rect 1026 1483 1037 1486
rect 1026 1416 1029 1476
rect 1018 1413 1029 1416
rect 986 1353 1005 1356
rect 978 1313 981 1336
rect 970 1243 981 1246
rect 978 1203 981 1243
rect 962 1123 965 1196
rect 962 863 965 1066
rect 970 1033 973 1196
rect 986 1156 989 1353
rect 994 1293 997 1346
rect 1010 1336 1013 1366
rect 1002 1333 1013 1336
rect 1002 1263 1005 1333
rect 1010 1313 1013 1326
rect 994 1213 997 1246
rect 1002 1203 1005 1226
rect 986 1153 997 1156
rect 970 983 973 1016
rect 970 903 973 936
rect 978 933 981 1136
rect 978 913 981 926
rect 962 803 965 826
rect 962 696 965 726
rect 970 703 973 896
rect 978 776 981 896
rect 986 783 989 1126
rect 994 1113 997 1153
rect 1002 1106 1005 1196
rect 994 1103 1005 1106
rect 994 876 997 1103
rect 1002 893 1005 1096
rect 1010 1083 1013 1216
rect 1018 1183 1021 1413
rect 1018 1133 1021 1176
rect 1018 1076 1021 1106
rect 1010 1073 1021 1076
rect 1010 1013 1013 1073
rect 1018 993 1021 1026
rect 1010 913 1013 986
rect 1018 913 1021 936
rect 1018 893 1021 906
rect 994 873 1001 876
rect 998 816 1001 873
rect 998 813 1005 816
rect 978 773 989 776
rect 962 693 973 696
rect 906 463 917 466
rect 930 513 941 516
rect 874 413 885 416
rect 890 393 893 406
rect 874 323 885 326
rect 858 293 869 296
rect 858 246 861 293
rect 874 263 877 316
rect 858 243 869 246
rect 866 226 869 243
rect 866 223 885 226
rect 874 196 877 216
rect 866 193 877 196
rect 834 123 837 156
rect 842 133 845 186
rect 858 133 861 146
rect 866 133 869 166
rect 786 93 797 96
rect 786 73 789 93
rect 850 43 853 126
rect 882 123 885 223
rect 890 193 893 316
rect 898 63 901 416
rect 906 413 909 463
rect 930 403 933 513
rect 906 333 909 356
rect 906 203 909 316
rect 914 303 917 326
rect 914 183 917 216
rect 922 213 925 226
rect 938 203 941 496
rect 946 433 949 656
rect 954 613 965 616
rect 954 603 965 606
rect 970 603 973 693
rect 978 683 981 736
rect 986 716 989 773
rect 994 723 997 756
rect 1002 733 1005 813
rect 986 713 997 716
rect 978 596 981 606
rect 962 593 981 596
rect 954 513 957 566
rect 962 523 965 593
rect 986 583 989 706
rect 994 573 997 713
rect 1002 683 1005 726
rect 1010 686 1013 866
rect 1018 823 1021 846
rect 1018 703 1021 796
rect 1010 683 1017 686
rect 962 506 965 516
rect 978 513 981 526
rect 994 513 997 526
rect 962 503 973 506
rect 970 446 973 503
rect 986 496 989 506
rect 1002 503 1005 676
rect 1014 536 1017 683
rect 1010 533 1017 536
rect 986 493 1005 496
rect 962 443 973 446
rect 962 356 965 443
rect 978 376 981 436
rect 986 396 989 476
rect 994 403 997 436
rect 1002 413 1005 446
rect 1002 396 1005 406
rect 986 393 1005 396
rect 978 373 989 376
rect 986 356 989 373
rect 962 353 973 356
rect 954 333 965 336
rect 954 303 957 326
rect 970 323 973 353
rect 978 333 981 356
rect 986 353 993 356
rect 978 296 981 326
rect 970 293 981 296
rect 990 286 993 353
rect 1002 313 1005 393
rect 1010 333 1013 533
rect 1018 373 1021 516
rect 1026 393 1029 1406
rect 1034 623 1037 1483
rect 1050 1446 1053 1563
rect 1062 1526 1065 1603
rect 1074 1583 1077 1603
rect 1074 1533 1077 1556
rect 1062 1523 1069 1526
rect 1042 1443 1053 1446
rect 1042 1383 1045 1443
rect 1042 1313 1045 1376
rect 1042 1093 1045 1296
rect 1050 1233 1053 1416
rect 1058 1326 1061 1426
rect 1066 1376 1069 1523
rect 1082 1523 1093 1526
rect 1082 1506 1085 1523
rect 1078 1503 1085 1506
rect 1078 1426 1081 1503
rect 1078 1423 1085 1426
rect 1074 1383 1077 1406
rect 1082 1403 1085 1423
rect 1066 1373 1077 1376
rect 1066 1333 1069 1373
rect 1058 1323 1069 1326
rect 1042 1063 1045 1086
rect 1050 1053 1053 1226
rect 1058 1193 1061 1316
rect 1058 1133 1061 1186
rect 1050 1013 1053 1026
rect 1042 896 1045 1006
rect 1058 1003 1061 1126
rect 1066 1023 1069 1323
rect 1074 1313 1077 1326
rect 1050 913 1053 996
rect 1058 943 1061 986
rect 1066 943 1069 996
rect 1058 903 1061 936
rect 1042 893 1049 896
rect 1046 796 1049 893
rect 1058 803 1061 826
rect 1066 813 1069 866
rect 1074 846 1077 1266
rect 1082 1193 1085 1366
rect 1082 863 1085 1136
rect 1074 843 1085 846
rect 1074 806 1077 836
rect 1066 803 1077 806
rect 1046 793 1077 796
rect 1034 413 1037 616
rect 1042 603 1045 736
rect 1026 356 1029 386
rect 1022 353 1029 356
rect 1022 296 1025 353
rect 1042 336 1045 576
rect 1050 456 1053 786
rect 1058 603 1061 746
rect 1066 623 1069 786
rect 1074 706 1077 793
rect 1082 723 1085 843
rect 1074 703 1081 706
rect 1066 596 1069 616
rect 1058 593 1069 596
rect 1058 513 1061 593
rect 1078 586 1081 703
rect 1090 613 1093 1516
rect 1098 1503 1101 1783
rect 1098 1363 1101 1416
rect 1098 1223 1101 1336
rect 1098 1136 1101 1156
rect 1106 1146 1109 1626
rect 1114 1403 1117 1863
rect 1154 1836 1157 1916
rect 1162 1893 1165 2006
rect 1122 1803 1125 1836
rect 1146 1833 1157 1836
rect 1130 1723 1141 1726
rect 1130 1693 1133 1716
rect 1138 1703 1141 1716
rect 1122 1623 1125 1676
rect 1122 1513 1125 1546
rect 1122 1413 1125 1426
rect 1114 1323 1117 1366
rect 1122 1293 1125 1406
rect 1130 1383 1133 1666
rect 1146 1646 1149 1833
rect 1154 1823 1165 1826
rect 1154 1733 1157 1756
rect 1146 1643 1157 1646
rect 1146 1623 1149 1636
rect 1138 1523 1141 1616
rect 1146 1416 1149 1536
rect 1154 1473 1157 1643
rect 1146 1413 1153 1416
rect 1130 1303 1133 1376
rect 1114 1223 1117 1246
rect 1122 1213 1125 1276
rect 1114 1173 1117 1206
rect 1130 1203 1133 1246
rect 1138 1226 1141 1406
rect 1150 1346 1153 1413
rect 1162 1403 1165 1816
rect 1170 1663 1173 2033
rect 1178 2003 1181 2196
rect 1186 2133 1189 2146
rect 1178 1933 1181 1986
rect 1186 1913 1189 2106
rect 1194 1943 1197 2203
rect 1206 2146 1209 2213
rect 1206 2143 1213 2146
rect 1218 2143 1221 2206
rect 1242 2156 1245 2216
rect 1258 2203 1261 2223
rect 1266 2186 1269 2276
rect 1250 2183 1269 2186
rect 1250 2173 1253 2183
rect 1234 2153 1245 2156
rect 1202 2123 1205 2136
rect 1210 2133 1213 2143
rect 1202 1976 1205 2026
rect 1210 1986 1213 2016
rect 1218 1996 1221 2056
rect 1226 2003 1229 2036
rect 1218 1993 1229 1996
rect 1210 1983 1229 1986
rect 1202 1973 1221 1976
rect 1178 1813 1181 1826
rect 1186 1803 1189 1856
rect 1210 1826 1213 1936
rect 1218 1923 1221 1973
rect 1226 1933 1229 1983
rect 1234 1953 1237 2153
rect 1242 2143 1253 2146
rect 1258 2096 1261 2166
rect 1266 2133 1269 2176
rect 1274 2123 1277 2226
rect 1274 2096 1277 2116
rect 1258 2093 1277 2096
rect 1242 1946 1245 2006
rect 1258 2003 1261 2016
rect 1234 1943 1245 1946
rect 1250 1976 1253 1996
rect 1266 1993 1269 2086
rect 1282 2076 1285 2476
rect 1290 2473 1301 2476
rect 1322 2483 1333 2486
rect 1338 2483 1345 2486
rect 1290 2396 1293 2473
rect 1298 2403 1301 2446
rect 1306 2403 1309 2436
rect 1314 2413 1317 2426
rect 1290 2393 1301 2396
rect 1290 2306 1293 2386
rect 1298 2323 1301 2393
rect 1322 2346 1325 2483
rect 1338 2463 1341 2483
rect 1354 2456 1357 2573
rect 1386 2546 1389 2616
rect 1410 2613 1413 2736
rect 1434 2686 1437 2726
rect 1430 2683 1437 2686
rect 1430 2606 1433 2683
rect 1446 2676 1449 2743
rect 1442 2673 1449 2676
rect 1442 2613 1445 2673
rect 1430 2603 1437 2606
rect 1434 2556 1437 2603
rect 1458 2586 1461 2776
rect 1558 2766 1561 2843
rect 1570 2813 1573 2936
rect 1594 2933 1597 3036
rect 1610 3026 1613 3116
rect 1650 3096 1653 3116
rect 1658 3113 1669 3116
rect 1642 3093 1653 3096
rect 1642 3046 1645 3093
rect 1642 3043 1653 3046
rect 1610 3023 1629 3026
rect 1650 3023 1653 3043
rect 1666 3036 1669 3113
rect 1714 3096 1717 3116
rect 1706 3093 1717 3096
rect 1722 3096 1725 3116
rect 1754 3106 1757 3136
rect 1738 3103 1757 3106
rect 1722 3093 1729 3096
rect 1706 3046 1709 3093
rect 1706 3043 1717 3046
rect 1658 3033 1669 3036
rect 1618 2976 1621 3016
rect 1626 3006 1629 3023
rect 1634 3013 1645 3016
rect 1626 3003 1653 3006
rect 1602 2973 1621 2976
rect 1602 2926 1605 2973
rect 1658 2966 1661 3033
rect 1714 3026 1717 3043
rect 1726 3036 1729 3093
rect 1726 3033 1733 3036
rect 1714 3023 1725 3026
rect 1674 3013 1693 3016
rect 1666 2973 1669 2996
rect 1594 2923 1605 2926
rect 1618 2963 1661 2966
rect 1618 2923 1621 2963
rect 1658 2933 1661 2946
rect 1554 2763 1561 2766
rect 1482 2723 1493 2726
rect 1514 2676 1517 2736
rect 1474 2673 1517 2676
rect 1474 2603 1477 2673
rect 1538 2626 1541 2726
rect 1554 2676 1557 2763
rect 1578 2726 1581 2816
rect 1594 2813 1597 2923
rect 1650 2886 1653 2926
rect 1658 2903 1661 2926
rect 1618 2883 1653 2886
rect 1618 2813 1621 2883
rect 1586 2793 1589 2806
rect 1594 2803 1605 2806
rect 1626 2763 1629 2816
rect 1634 2783 1637 2806
rect 1642 2746 1645 2856
rect 1658 2813 1661 2886
rect 1674 2853 1677 3013
rect 1682 2933 1685 2966
rect 1690 2913 1693 3006
rect 1706 3003 1709 3016
rect 1722 2946 1725 3023
rect 1730 3003 1733 3033
rect 1730 2973 1733 2996
rect 1722 2943 1733 2946
rect 1706 2886 1709 2936
rect 1698 2883 1709 2886
rect 1698 2836 1701 2883
rect 1730 2856 1733 2943
rect 1738 2923 1741 3103
rect 1762 3096 1765 3136
rect 1746 3093 1765 3096
rect 1778 3133 1789 3136
rect 1802 3136 1805 3166
rect 1810 3146 1813 3216
rect 1810 3143 1845 3146
rect 1802 3133 1821 3136
rect 1842 3133 1845 3143
rect 1850 3133 1853 3146
rect 1746 3003 1749 3093
rect 1778 3076 1781 3133
rect 1794 3083 1797 3126
rect 1810 3123 1813 3133
rect 1874 3126 1877 3216
rect 1890 3183 1893 3206
rect 1938 3176 1941 3216
rect 1938 3173 1973 3176
rect 1818 3116 1821 3126
rect 1826 3123 1877 3126
rect 1802 3113 1813 3116
rect 1818 3113 1845 3116
rect 1778 3073 1821 3076
rect 1754 3013 1757 3026
rect 1762 3013 1765 3046
rect 1754 2993 1757 3006
rect 1770 2966 1773 3026
rect 1778 3003 1781 3016
rect 1786 3013 1797 3016
rect 1802 3013 1805 3066
rect 1818 3056 1821 3073
rect 1818 3053 1825 3056
rect 1794 2983 1797 3006
rect 1802 2993 1805 3006
rect 1770 2963 1777 2966
rect 1774 2886 1777 2963
rect 1722 2853 1733 2856
rect 1770 2883 1777 2886
rect 1786 2883 1789 2926
rect 1810 2903 1813 3026
rect 1822 2996 1825 3053
rect 1834 3003 1845 3006
rect 1822 2993 1837 2996
rect 1650 2753 1653 2806
rect 1666 2783 1669 2816
rect 1674 2766 1677 2836
rect 1698 2833 1709 2836
rect 1722 2833 1725 2853
rect 1706 2813 1709 2833
rect 1770 2823 1773 2883
rect 1682 2793 1685 2806
rect 1670 2763 1677 2766
rect 1642 2743 1653 2746
rect 1578 2723 1597 2726
rect 1626 2723 1629 2736
rect 1554 2673 1565 2676
rect 1562 2656 1565 2673
rect 1562 2653 1573 2656
rect 1530 2623 1541 2626
rect 1458 2583 1477 2586
rect 1346 2453 1357 2456
rect 1370 2543 1389 2546
rect 1402 2553 1437 2556
rect 1338 2356 1341 2426
rect 1346 2413 1349 2453
rect 1306 2343 1325 2346
rect 1334 2353 1341 2356
rect 1290 2303 1297 2306
rect 1294 2236 1297 2303
rect 1278 2073 1285 2076
rect 1290 2233 1297 2236
rect 1278 2016 1281 2073
rect 1290 2033 1293 2233
rect 1298 2016 1301 2216
rect 1306 2026 1309 2343
rect 1314 2303 1317 2336
rect 1314 2223 1317 2286
rect 1314 2113 1317 2126
rect 1306 2023 1317 2026
rect 1278 2013 1285 2016
rect 1250 1973 1261 1976
rect 1234 1836 1237 1943
rect 1242 1923 1245 1936
rect 1250 1933 1253 1973
rect 1250 1913 1253 1926
rect 1234 1833 1245 1836
rect 1210 1823 1229 1826
rect 1210 1803 1213 1816
rect 1178 1723 1181 1736
rect 1178 1636 1181 1646
rect 1170 1633 1181 1636
rect 1170 1423 1173 1536
rect 1178 1533 1181 1546
rect 1186 1533 1189 1716
rect 1218 1713 1221 1736
rect 1226 1696 1229 1823
rect 1234 1786 1237 1816
rect 1242 1803 1245 1833
rect 1258 1816 1261 1966
rect 1266 1916 1269 1946
rect 1274 1923 1277 1996
rect 1266 1913 1273 1916
rect 1270 1826 1273 1913
rect 1270 1823 1277 1826
rect 1254 1813 1261 1816
rect 1234 1783 1245 1786
rect 1242 1736 1245 1783
rect 1254 1756 1257 1813
rect 1274 1806 1277 1823
rect 1282 1813 1285 2013
rect 1290 2003 1293 2016
rect 1298 2013 1317 2016
rect 1290 1953 1293 1996
rect 1298 1963 1301 2006
rect 1290 1926 1293 1946
rect 1290 1923 1297 1926
rect 1306 1923 1309 2006
rect 1294 1846 1297 1923
rect 1306 1863 1309 1916
rect 1314 1846 1317 2013
rect 1290 1843 1297 1846
rect 1310 1843 1317 1846
rect 1254 1753 1261 1756
rect 1234 1733 1245 1736
rect 1258 1733 1261 1753
rect 1234 1713 1237 1733
rect 1266 1716 1269 1806
rect 1274 1803 1285 1806
rect 1258 1713 1269 1716
rect 1194 1516 1197 1626
rect 1202 1593 1205 1606
rect 1190 1513 1197 1516
rect 1178 1416 1181 1466
rect 1190 1436 1193 1513
rect 1190 1433 1197 1436
rect 1170 1413 1181 1416
rect 1178 1393 1181 1406
rect 1146 1343 1153 1346
rect 1146 1236 1149 1343
rect 1162 1326 1165 1336
rect 1154 1323 1165 1326
rect 1154 1243 1157 1323
rect 1162 1293 1165 1316
rect 1146 1233 1157 1236
rect 1138 1223 1149 1226
rect 1122 1166 1125 1186
rect 1122 1163 1133 1166
rect 1106 1143 1125 1146
rect 1098 1133 1109 1136
rect 1098 1123 1109 1126
rect 1114 1103 1117 1126
rect 1122 1096 1125 1143
rect 1130 1133 1133 1163
rect 1138 1133 1141 1216
rect 1146 1193 1149 1223
rect 1154 1146 1157 1233
rect 1146 1143 1157 1146
rect 1098 1023 1101 1096
rect 1106 1093 1125 1096
rect 1098 933 1101 1016
rect 1106 926 1109 1093
rect 1114 946 1117 1066
rect 1122 1013 1125 1026
rect 1130 1023 1133 1086
rect 1138 1063 1141 1116
rect 1122 953 1125 986
rect 1130 953 1133 966
rect 1114 943 1133 946
rect 1098 923 1109 926
rect 1114 923 1117 936
rect 1130 916 1133 943
rect 1114 913 1133 916
rect 1098 733 1101 826
rect 1098 693 1101 726
rect 1106 676 1109 906
rect 1114 813 1117 913
rect 1114 783 1117 806
rect 1102 673 1109 676
rect 1102 606 1105 673
rect 1114 653 1117 736
rect 1114 613 1117 646
rect 1122 613 1125 906
rect 1130 886 1133 906
rect 1138 893 1141 1016
rect 1146 896 1149 1143
rect 1162 1136 1165 1226
rect 1154 1133 1165 1136
rect 1170 1136 1173 1386
rect 1186 1376 1189 1416
rect 1182 1373 1189 1376
rect 1182 1316 1185 1373
rect 1178 1313 1185 1316
rect 1178 1153 1181 1313
rect 1194 1306 1197 1433
rect 1186 1303 1197 1306
rect 1186 1243 1189 1303
rect 1170 1133 1177 1136
rect 1154 903 1157 1133
rect 1162 1003 1165 1126
rect 1174 1026 1177 1133
rect 1186 1063 1189 1216
rect 1194 1203 1197 1296
rect 1194 1133 1197 1196
rect 1170 1023 1177 1026
rect 1194 1023 1197 1086
rect 1170 996 1173 1023
rect 1162 993 1173 996
rect 1178 1003 1189 1006
rect 1162 916 1165 993
rect 1178 926 1181 1003
rect 1170 923 1181 926
rect 1186 923 1189 966
rect 1194 916 1197 1006
rect 1162 913 1173 916
rect 1146 893 1165 896
rect 1130 883 1149 886
rect 1130 823 1133 866
rect 1130 793 1133 806
rect 1138 733 1141 836
rect 1146 726 1149 883
rect 1154 753 1157 826
rect 1162 746 1165 893
rect 1170 796 1173 913
rect 1178 803 1181 916
rect 1186 913 1197 916
rect 1186 813 1189 913
rect 1194 843 1197 896
rect 1202 796 1205 1586
rect 1210 903 1213 1696
rect 1226 1693 1233 1696
rect 1218 1613 1221 1666
rect 1230 1626 1233 1693
rect 1258 1646 1261 1713
rect 1258 1643 1269 1646
rect 1226 1623 1233 1626
rect 1226 1606 1229 1623
rect 1242 1613 1245 1626
rect 1218 1603 1229 1606
rect 1218 1466 1221 1603
rect 1250 1556 1253 1606
rect 1258 1573 1261 1616
rect 1226 1483 1229 1556
rect 1234 1553 1253 1556
rect 1218 1463 1225 1466
rect 1222 1386 1225 1463
rect 1218 1383 1225 1386
rect 1218 1363 1221 1383
rect 1218 1303 1221 1336
rect 1218 1216 1221 1236
rect 1226 1223 1229 1336
rect 1218 1213 1229 1216
rect 1234 1196 1237 1553
rect 1242 1543 1261 1546
rect 1242 1523 1245 1543
rect 1250 1526 1253 1536
rect 1258 1533 1261 1543
rect 1266 1526 1269 1643
rect 1250 1523 1269 1526
rect 1250 1456 1253 1523
rect 1242 1453 1253 1456
rect 1242 1293 1245 1453
rect 1266 1423 1269 1496
rect 1250 1403 1253 1416
rect 1258 1393 1261 1416
rect 1250 1303 1253 1326
rect 1258 1286 1261 1336
rect 1242 1203 1245 1286
rect 1254 1283 1261 1286
rect 1254 1216 1257 1283
rect 1254 1213 1261 1216
rect 1234 1193 1253 1196
rect 1218 1123 1221 1136
rect 1250 1133 1253 1193
rect 1218 1103 1221 1116
rect 1242 1103 1245 1126
rect 1258 1116 1261 1213
rect 1266 1133 1269 1416
rect 1274 1403 1277 1736
rect 1282 1716 1285 1803
rect 1290 1723 1293 1843
rect 1282 1713 1289 1716
rect 1286 1656 1289 1713
rect 1286 1653 1293 1656
rect 1282 1523 1285 1636
rect 1290 1506 1293 1653
rect 1298 1623 1301 1826
rect 1310 1756 1313 1843
rect 1310 1753 1317 1756
rect 1314 1733 1317 1753
rect 1322 1723 1325 2316
rect 1334 2306 1337 2353
rect 1354 2333 1357 2416
rect 1362 2393 1365 2436
rect 1370 2403 1373 2543
rect 1386 2523 1389 2536
rect 1394 2523 1397 2536
rect 1402 2496 1405 2553
rect 1410 2503 1413 2536
rect 1418 2523 1421 2546
rect 1426 2543 1461 2546
rect 1466 2543 1469 2576
rect 1426 2533 1429 2543
rect 1450 2526 1453 2536
rect 1458 2533 1461 2543
rect 1442 2523 1453 2526
rect 1442 2516 1445 2523
rect 1418 2513 1445 2516
rect 1458 2503 1461 2516
rect 1474 2496 1477 2583
rect 1482 2543 1485 2586
rect 1402 2493 1437 2496
rect 1394 2426 1397 2446
rect 1390 2423 1397 2426
rect 1378 2346 1381 2416
rect 1390 2376 1393 2423
rect 1402 2386 1405 2436
rect 1410 2393 1413 2426
rect 1418 2413 1421 2426
rect 1426 2413 1429 2466
rect 1434 2416 1437 2493
rect 1458 2493 1477 2496
rect 1442 2423 1445 2446
rect 1458 2416 1461 2493
rect 1434 2413 1445 2416
rect 1450 2413 1461 2416
rect 1418 2396 1421 2406
rect 1442 2403 1445 2413
rect 1466 2396 1469 2466
rect 1418 2393 1429 2396
rect 1462 2393 1469 2396
rect 1418 2386 1421 2393
rect 1402 2383 1421 2386
rect 1390 2373 1397 2376
rect 1378 2343 1385 2346
rect 1334 2303 1341 2306
rect 1330 2213 1333 2246
rect 1338 2236 1341 2303
rect 1382 2296 1385 2343
rect 1378 2293 1385 2296
rect 1338 2233 1349 2236
rect 1338 2206 1341 2226
rect 1330 2203 1341 2206
rect 1330 2106 1333 2136
rect 1338 2123 1341 2196
rect 1330 2103 1337 2106
rect 1334 2036 1337 2103
rect 1330 2033 1337 2036
rect 1330 1993 1333 2033
rect 1338 2003 1341 2016
rect 1346 1966 1349 2233
rect 1354 2143 1357 2246
rect 1362 2083 1365 2136
rect 1354 1983 1357 2006
rect 1330 1953 1333 1966
rect 1338 1963 1349 1966
rect 1338 1946 1341 1963
rect 1354 1946 1357 1966
rect 1330 1943 1341 1946
rect 1350 1943 1357 1946
rect 1362 1943 1365 2036
rect 1370 2013 1373 2186
rect 1378 2116 1381 2293
rect 1386 2203 1389 2226
rect 1386 2133 1389 2146
rect 1378 2113 1385 2116
rect 1382 2026 1385 2113
rect 1394 2093 1397 2373
rect 1402 2303 1405 2326
rect 1426 2316 1429 2376
rect 1434 2323 1437 2336
rect 1442 2323 1445 2386
rect 1450 2333 1453 2356
rect 1426 2313 1437 2316
rect 1402 2233 1421 2236
rect 1402 2133 1405 2186
rect 1410 2116 1413 2226
rect 1418 2203 1421 2233
rect 1406 2113 1413 2116
rect 1406 2026 1409 2113
rect 1378 2023 1385 2026
rect 1378 1996 1381 2023
rect 1394 2013 1397 2026
rect 1406 2023 1413 2026
rect 1374 1993 1381 1996
rect 1306 1673 1309 1716
rect 1330 1686 1333 1943
rect 1338 1903 1341 1936
rect 1338 1813 1341 1886
rect 1350 1876 1353 1943
rect 1350 1873 1357 1876
rect 1338 1763 1341 1806
rect 1346 1803 1349 1856
rect 1354 1786 1357 1873
rect 1362 1863 1365 1936
rect 1374 1906 1377 1993
rect 1386 1933 1389 2006
rect 1374 1903 1381 1906
rect 1378 1883 1381 1903
rect 1386 1866 1389 1916
rect 1382 1863 1389 1866
rect 1350 1783 1357 1786
rect 1362 1823 1373 1826
rect 1322 1683 1333 1686
rect 1322 1636 1325 1683
rect 1322 1633 1329 1636
rect 1286 1503 1293 1506
rect 1286 1436 1289 1503
rect 1282 1433 1289 1436
rect 1282 1383 1285 1433
rect 1274 1263 1277 1326
rect 1282 1313 1285 1346
rect 1282 1186 1285 1216
rect 1290 1203 1293 1426
rect 1298 1423 1301 1606
rect 1298 1323 1301 1386
rect 1254 1113 1261 1116
rect 1218 926 1221 1026
rect 1226 936 1229 1066
rect 1254 1036 1257 1113
rect 1254 1033 1261 1036
rect 1234 1003 1237 1026
rect 1242 1013 1253 1016
rect 1258 996 1261 1033
rect 1250 993 1261 996
rect 1226 933 1237 936
rect 1218 923 1229 926
rect 1170 793 1181 796
rect 1138 723 1149 726
rect 1154 743 1165 746
rect 1074 583 1081 586
rect 1090 603 1105 606
rect 1050 453 1069 456
rect 1058 366 1061 406
rect 1066 383 1069 453
rect 1058 363 1069 366
rect 1034 333 1045 336
rect 1034 306 1037 326
rect 1066 323 1069 363
rect 1074 333 1077 583
rect 1082 503 1085 516
rect 1090 446 1093 603
rect 1098 566 1101 586
rect 1098 563 1105 566
rect 1102 486 1105 563
rect 1114 503 1117 606
rect 1102 483 1109 486
rect 1090 443 1097 446
rect 1082 423 1085 436
rect 1094 396 1097 443
rect 1090 393 1097 396
rect 1082 333 1085 376
rect 1034 303 1045 306
rect 986 283 993 286
rect 1018 293 1025 296
rect 962 193 965 226
rect 986 183 989 283
rect 1018 226 1021 293
rect 1042 246 1045 303
rect 1090 276 1093 393
rect 1106 376 1109 483
rect 1130 426 1133 696
rect 1138 616 1141 723
rect 1154 706 1157 743
rect 1150 703 1157 706
rect 1150 636 1153 703
rect 1150 633 1157 636
rect 1138 613 1149 616
rect 1154 596 1157 633
rect 1150 593 1157 596
rect 1138 503 1141 526
rect 1150 496 1153 593
rect 1162 503 1165 726
rect 1170 556 1173 656
rect 1178 573 1181 793
rect 1194 793 1205 796
rect 1194 696 1197 793
rect 1194 693 1205 696
rect 1186 603 1189 616
rect 1194 613 1197 676
rect 1170 553 1177 556
rect 1174 496 1177 553
rect 1150 493 1157 496
rect 1130 423 1141 426
rect 1034 243 1045 246
rect 1082 273 1093 276
rect 1098 373 1109 376
rect 1122 373 1125 406
rect 1034 226 1037 243
rect 1082 226 1085 273
rect 1098 226 1101 373
rect 1114 323 1117 356
rect 1106 303 1109 316
rect 1122 306 1125 336
rect 1118 303 1125 306
rect 1106 233 1109 256
rect 1018 223 1029 226
rect 1034 223 1053 226
rect 1082 223 1093 226
rect 1098 223 1109 226
rect 1026 203 1029 223
rect 1034 213 1053 216
rect 1050 146 1053 206
rect 1090 203 1093 223
rect 1118 206 1121 303
rect 1114 203 1121 206
rect 946 143 973 146
rect 938 93 941 136
rect 946 123 949 143
rect 970 133 973 143
rect 1034 143 1053 146
rect 1026 116 1029 126
rect 1034 123 1037 143
rect 1066 133 1069 156
rect 1114 146 1117 203
rect 1114 143 1125 146
rect 1122 126 1125 143
rect 1130 133 1133 326
rect 1138 306 1141 423
rect 1146 406 1149 476
rect 1154 413 1157 493
rect 1170 493 1177 496
rect 1170 413 1173 493
rect 1186 486 1189 536
rect 1194 523 1197 606
rect 1202 543 1205 693
rect 1202 503 1205 526
rect 1210 513 1213 856
rect 1218 823 1221 866
rect 1218 486 1221 756
rect 1226 653 1229 923
rect 1234 903 1237 926
rect 1242 913 1245 936
rect 1250 906 1253 993
rect 1266 976 1269 1086
rect 1274 1023 1277 1186
rect 1282 1183 1289 1186
rect 1286 1026 1289 1183
rect 1282 1023 1289 1026
rect 1282 986 1285 1023
rect 1298 1013 1301 1256
rect 1306 1236 1309 1606
rect 1314 1523 1317 1616
rect 1326 1566 1329 1633
rect 1326 1563 1333 1566
rect 1330 1543 1333 1563
rect 1314 1343 1317 1486
rect 1322 1326 1325 1516
rect 1330 1343 1333 1456
rect 1314 1323 1325 1326
rect 1314 1253 1317 1323
rect 1322 1293 1325 1316
rect 1306 1233 1313 1236
rect 1310 1146 1313 1233
rect 1322 1173 1325 1256
rect 1330 1183 1333 1336
rect 1306 1143 1313 1146
rect 1262 973 1269 976
rect 1274 983 1285 986
rect 1262 916 1265 973
rect 1274 933 1277 983
rect 1262 913 1269 916
rect 1242 903 1253 906
rect 1242 876 1245 903
rect 1250 893 1261 896
rect 1250 883 1253 893
rect 1266 876 1269 913
rect 1234 873 1245 876
rect 1262 873 1269 876
rect 1234 853 1237 873
rect 1234 706 1237 806
rect 1242 726 1245 866
rect 1250 813 1253 836
rect 1262 796 1265 873
rect 1274 863 1277 926
rect 1274 803 1277 846
rect 1282 833 1285 976
rect 1282 803 1285 816
rect 1262 793 1269 796
rect 1250 733 1253 786
rect 1242 723 1253 726
rect 1234 703 1241 706
rect 1238 646 1241 703
rect 1234 643 1241 646
rect 1234 623 1237 643
rect 1226 583 1229 616
rect 1186 483 1197 486
rect 1194 406 1197 483
rect 1146 403 1157 406
rect 1146 323 1149 336
rect 1138 303 1145 306
rect 1142 156 1145 303
rect 1154 186 1157 403
rect 1162 386 1165 406
rect 1186 403 1197 406
rect 1210 483 1221 486
rect 1162 383 1169 386
rect 1166 326 1169 383
rect 1186 336 1189 403
rect 1210 346 1213 483
rect 1226 416 1229 516
rect 1242 513 1245 526
rect 1250 503 1253 723
rect 1266 693 1269 793
rect 1274 723 1277 736
rect 1290 626 1293 1006
rect 1298 943 1301 986
rect 1298 813 1301 936
rect 1298 783 1301 806
rect 1306 736 1309 1143
rect 1322 1133 1325 1146
rect 1314 1106 1317 1126
rect 1314 1103 1321 1106
rect 1318 1036 1321 1103
rect 1318 1033 1325 1036
rect 1314 1003 1317 1016
rect 1322 1003 1325 1033
rect 1314 763 1317 936
rect 1322 766 1325 996
rect 1330 773 1333 1156
rect 1338 1043 1341 1676
rect 1350 1666 1353 1783
rect 1350 1663 1357 1666
rect 1346 1623 1349 1646
rect 1346 1553 1349 1616
rect 1346 1533 1349 1546
rect 1354 1516 1357 1663
rect 1362 1586 1365 1823
rect 1370 1803 1373 1816
rect 1382 1746 1385 1863
rect 1370 1723 1373 1746
rect 1382 1743 1389 1746
rect 1378 1713 1381 1726
rect 1370 1603 1373 1706
rect 1386 1696 1389 1743
rect 1394 1733 1397 1926
rect 1402 1903 1405 2006
rect 1410 1976 1413 2023
rect 1418 1986 1421 2186
rect 1426 1996 1429 2206
rect 1434 2193 1437 2313
rect 1462 2306 1465 2393
rect 1474 2356 1477 2416
rect 1490 2413 1493 2526
rect 1498 2483 1501 2606
rect 1530 2566 1533 2623
rect 1530 2563 1541 2566
rect 1506 2523 1509 2536
rect 1514 2523 1517 2556
rect 1522 2516 1525 2536
rect 1530 2533 1533 2546
rect 1538 2536 1541 2563
rect 1546 2546 1549 2616
rect 1570 2596 1573 2653
rect 1562 2593 1573 2596
rect 1562 2573 1565 2593
rect 1546 2543 1589 2546
rect 1538 2533 1549 2536
rect 1522 2513 1533 2516
rect 1506 2403 1509 2456
rect 1530 2413 1533 2513
rect 1538 2483 1541 2526
rect 1546 2423 1549 2533
rect 1554 2533 1565 2536
rect 1554 2523 1557 2533
rect 1562 2516 1565 2526
rect 1570 2523 1573 2536
rect 1586 2533 1589 2543
rect 1594 2533 1597 2546
rect 1602 2543 1605 2566
rect 1554 2503 1557 2516
rect 1562 2513 1589 2516
rect 1610 2463 1613 2626
rect 1618 2543 1621 2616
rect 1626 2543 1629 2596
rect 1642 2546 1645 2616
rect 1634 2543 1645 2546
rect 1634 2473 1637 2543
rect 1650 2536 1653 2743
rect 1658 2623 1661 2726
rect 1670 2686 1673 2763
rect 1690 2706 1693 2746
rect 1706 2723 1709 2766
rect 1722 2743 1725 2806
rect 1690 2703 1701 2706
rect 1738 2703 1741 2726
rect 1670 2683 1677 2686
rect 1658 2593 1661 2616
rect 1674 2553 1677 2683
rect 1698 2646 1701 2703
rect 1690 2643 1701 2646
rect 1690 2596 1693 2643
rect 1698 2603 1701 2616
rect 1690 2593 1701 2596
rect 1642 2533 1653 2536
rect 1658 2533 1677 2536
rect 1682 2533 1685 2546
rect 1690 2543 1693 2566
rect 1594 2423 1637 2426
rect 1594 2413 1597 2423
rect 1474 2353 1517 2356
rect 1458 2303 1465 2306
rect 1474 2303 1477 2336
rect 1458 2236 1461 2303
rect 1458 2233 1469 2236
rect 1458 2146 1461 2216
rect 1434 2143 1461 2146
rect 1434 2013 1437 2143
rect 1442 2106 1445 2116
rect 1450 2106 1453 2116
rect 1442 2103 1453 2106
rect 1442 2043 1445 2103
rect 1442 2003 1445 2036
rect 1426 1993 1445 1996
rect 1418 1983 1429 1986
rect 1410 1973 1421 1976
rect 1410 1796 1413 1966
rect 1418 1873 1421 1973
rect 1426 1813 1429 1983
rect 1434 1876 1437 1936
rect 1442 1883 1445 1993
rect 1434 1873 1445 1876
rect 1434 1813 1437 1866
rect 1442 1813 1445 1873
rect 1418 1803 1429 1806
rect 1434 1803 1445 1806
rect 1410 1793 1421 1796
rect 1394 1713 1397 1726
rect 1386 1693 1393 1696
rect 1378 1603 1381 1666
rect 1390 1626 1393 1693
rect 1386 1623 1393 1626
rect 1386 1603 1389 1623
rect 1362 1583 1369 1586
rect 1350 1513 1357 1516
rect 1350 1436 1353 1513
rect 1366 1506 1369 1583
rect 1362 1503 1369 1506
rect 1362 1483 1365 1503
rect 1350 1433 1357 1436
rect 1346 1253 1349 1416
rect 1346 1223 1349 1236
rect 1338 993 1341 1006
rect 1346 986 1349 1176
rect 1338 983 1349 986
rect 1338 933 1341 983
rect 1346 923 1349 946
rect 1338 793 1341 866
rect 1322 763 1333 766
rect 1314 743 1317 756
rect 1330 743 1333 763
rect 1306 733 1325 736
rect 1338 733 1341 766
rect 1322 726 1325 733
rect 1274 623 1293 626
rect 1274 606 1277 623
rect 1282 613 1293 616
rect 1298 613 1309 616
rect 1266 596 1269 606
rect 1274 603 1285 606
rect 1290 603 1301 606
rect 1266 593 1277 596
rect 1274 543 1277 593
rect 1282 536 1285 603
rect 1266 533 1285 536
rect 1298 533 1301 603
rect 1222 413 1229 416
rect 1242 413 1245 426
rect 1258 413 1261 526
rect 1266 496 1269 533
rect 1306 526 1309 613
rect 1314 603 1317 726
rect 1322 723 1341 726
rect 1322 603 1325 646
rect 1298 523 1309 526
rect 1306 506 1309 523
rect 1298 503 1309 506
rect 1266 493 1285 496
rect 1222 366 1225 413
rect 1282 406 1285 493
rect 1222 363 1229 366
rect 1234 363 1237 406
rect 1250 373 1253 406
rect 1274 403 1285 406
rect 1210 343 1221 346
rect 1178 326 1181 336
rect 1186 333 1197 336
rect 1166 323 1189 326
rect 1194 316 1197 333
rect 1162 263 1165 316
rect 1186 313 1197 316
rect 1210 313 1213 326
rect 1170 283 1173 306
rect 1162 223 1165 256
rect 1186 236 1189 313
rect 1194 303 1213 306
rect 1178 233 1189 236
rect 1162 193 1165 216
rect 1154 183 1165 186
rect 1138 153 1145 156
rect 1042 123 1053 126
rect 1082 123 1125 126
rect 1042 116 1045 123
rect 954 33 957 116
rect 1018 83 1021 116
rect 1026 113 1045 116
rect 1066 113 1101 116
rect 1138 113 1141 153
rect 1146 93 1149 136
rect 1154 123 1157 166
rect 1162 136 1165 183
rect 1178 156 1181 233
rect 1194 206 1197 226
rect 1202 223 1205 256
rect 1194 203 1205 206
rect 1178 153 1189 156
rect 1162 133 1181 136
rect 1162 123 1173 126
rect 1162 83 1165 123
rect 1178 116 1181 133
rect 1186 123 1189 153
rect 1194 123 1197 203
rect 1210 196 1213 276
rect 1218 246 1221 343
rect 1226 263 1229 363
rect 1274 336 1277 403
rect 1298 396 1301 503
rect 1298 393 1309 396
rect 1306 373 1309 393
rect 1250 323 1253 336
rect 1266 333 1277 336
rect 1242 313 1253 316
rect 1218 243 1229 246
rect 1202 193 1213 196
rect 1202 116 1205 193
rect 1226 166 1229 243
rect 1250 233 1253 313
rect 1266 236 1269 333
rect 1314 316 1317 526
rect 1330 423 1333 616
rect 1338 596 1341 723
rect 1346 603 1349 616
rect 1338 593 1349 596
rect 1346 523 1349 593
rect 1338 416 1341 436
rect 1322 413 1341 416
rect 1322 403 1325 413
rect 1354 406 1357 1433
rect 1362 1413 1365 1456
rect 1378 1413 1381 1586
rect 1386 1453 1389 1516
rect 1362 1096 1365 1346
rect 1370 1133 1373 1406
rect 1378 1393 1381 1406
rect 1386 1373 1389 1416
rect 1378 1343 1389 1346
rect 1362 1093 1369 1096
rect 1366 1006 1369 1093
rect 1362 1003 1369 1006
rect 1362 983 1365 1003
rect 1378 983 1381 1336
rect 1394 1296 1397 1536
rect 1402 1526 1405 1716
rect 1410 1663 1413 1736
rect 1418 1733 1421 1793
rect 1426 1713 1429 1803
rect 1450 1796 1453 2096
rect 1458 2013 1461 2136
rect 1458 1903 1461 1936
rect 1466 1923 1469 2233
rect 1474 2193 1477 2246
rect 1474 2143 1477 2176
rect 1474 2033 1477 2136
rect 1482 2033 1485 2316
rect 1514 2293 1517 2353
rect 1562 2323 1565 2336
rect 1594 2323 1597 2406
rect 1602 2363 1605 2416
rect 1610 2413 1621 2416
rect 1634 2413 1637 2423
rect 1610 2383 1613 2406
rect 1618 2333 1621 2396
rect 1634 2393 1637 2406
rect 1642 2336 1645 2533
rect 1674 2526 1677 2533
rect 1650 2503 1653 2526
rect 1658 2513 1661 2526
rect 1674 2523 1685 2526
rect 1690 2516 1693 2536
rect 1682 2513 1693 2516
rect 1682 2493 1685 2513
rect 1650 2403 1653 2476
rect 1658 2396 1661 2466
rect 1690 2433 1693 2446
rect 1674 2403 1677 2426
rect 1698 2423 1701 2593
rect 1714 2573 1717 2606
rect 1746 2536 1749 2816
rect 1794 2813 1805 2816
rect 1754 2713 1757 2736
rect 1778 2733 1781 2776
rect 1810 2736 1813 2816
rect 1834 2776 1837 2993
rect 1850 2913 1853 3016
rect 1866 3013 1869 3076
rect 1858 2983 1861 3006
rect 1866 3003 1877 3006
rect 1882 3003 1885 3086
rect 1890 2993 1893 3016
rect 1898 2983 1901 3006
rect 1906 2966 1909 3136
rect 1914 3133 1917 3146
rect 1930 3133 1933 3146
rect 1946 3143 1965 3146
rect 1946 3133 1949 3143
rect 1930 3123 1949 3126
rect 1954 3123 1957 3136
rect 1922 3003 1925 3026
rect 1946 2976 1949 3076
rect 1858 2963 1909 2966
rect 1922 2973 1949 2976
rect 1858 2923 1861 2963
rect 1922 2943 1925 2973
rect 1954 2966 1957 3046
rect 1962 3013 1965 3143
rect 1970 3133 1973 3173
rect 1978 3143 1981 3216
rect 1994 3193 1997 3206
rect 1978 3123 1989 3126
rect 1994 3036 1997 3056
rect 1990 3033 1997 3036
rect 1938 2963 1957 2966
rect 1890 2933 1917 2936
rect 1842 2886 1845 2906
rect 1842 2883 1853 2886
rect 1850 2803 1853 2883
rect 1858 2813 1869 2816
rect 1858 2793 1861 2806
rect 1834 2773 1845 2776
rect 1802 2733 1813 2736
rect 1762 2723 1789 2726
rect 1810 2723 1813 2733
rect 1818 2706 1821 2756
rect 1810 2703 1821 2706
rect 1810 2626 1813 2703
rect 1802 2623 1813 2626
rect 1762 2576 1765 2616
rect 1762 2573 1773 2576
rect 1706 2483 1709 2536
rect 1722 2533 1749 2536
rect 1722 2466 1725 2533
rect 1762 2526 1765 2546
rect 1770 2533 1773 2573
rect 1778 2546 1781 2586
rect 1802 2566 1805 2623
rect 1802 2563 1813 2566
rect 1778 2543 1797 2546
rect 1746 2506 1749 2526
rect 1754 2513 1757 2526
rect 1762 2523 1773 2526
rect 1786 2523 1797 2526
rect 1770 2513 1773 2523
rect 1722 2463 1733 2466
rect 1714 2443 1725 2446
rect 1682 2413 1709 2416
rect 1698 2403 1709 2406
rect 1634 2333 1645 2336
rect 1650 2393 1661 2396
rect 1714 2396 1717 2416
rect 1722 2403 1725 2443
rect 1714 2393 1725 2396
rect 1650 2333 1653 2393
rect 1658 2333 1661 2356
rect 1714 2336 1717 2393
rect 1730 2376 1733 2463
rect 1738 2383 1741 2506
rect 1746 2503 1757 2506
rect 1746 2486 1749 2503
rect 1746 2483 1757 2486
rect 1754 2426 1757 2483
rect 1746 2423 1757 2426
rect 1746 2403 1749 2423
rect 1778 2403 1781 2436
rect 1802 2413 1805 2536
rect 1810 2496 1813 2563
rect 1818 2513 1821 2616
rect 1810 2493 1817 2496
rect 1814 2416 1817 2493
rect 1826 2433 1829 2746
rect 1834 2703 1837 2726
rect 1842 2713 1845 2773
rect 1850 2733 1853 2786
rect 1866 2763 1869 2813
rect 1858 2723 1861 2736
rect 1874 2683 1877 2826
rect 1882 2786 1885 2836
rect 1890 2813 1893 2926
rect 1890 2793 1893 2806
rect 1898 2803 1901 2816
rect 1906 2786 1909 2796
rect 1882 2783 1909 2786
rect 1898 2733 1901 2746
rect 1906 2733 1909 2783
rect 1914 2756 1917 2933
rect 1922 2896 1925 2926
rect 1930 2916 1933 2936
rect 1938 2923 1941 2963
rect 1962 2956 1965 2966
rect 1954 2953 1965 2956
rect 1990 2956 1993 3033
rect 2002 3026 2005 3126
rect 2010 3076 2013 3136
rect 2018 3133 2021 3156
rect 2042 3136 2045 3216
rect 2074 3153 2077 3216
rect 2090 3193 2093 3206
rect 2138 3193 2141 3216
rect 2170 3213 2189 3216
rect 2034 3113 2037 3136
rect 2042 3133 2061 3136
rect 2122 3133 2125 3146
rect 2138 3143 2149 3146
rect 2082 3123 2101 3126
rect 2082 3106 2085 3123
rect 2074 3103 2085 3106
rect 2010 3073 2045 3076
rect 2002 3023 2021 3026
rect 1990 2953 1997 2956
rect 1954 2923 1957 2953
rect 1962 2916 1965 2946
rect 1930 2913 1949 2916
rect 1946 2903 1949 2913
rect 1954 2913 1965 2916
rect 1970 2913 1973 2926
rect 1954 2896 1957 2913
rect 1978 2903 1981 2936
rect 1986 2923 1989 2936
rect 1994 2923 1997 2953
rect 1922 2893 1957 2896
rect 1930 2816 1933 2866
rect 2002 2856 2005 3016
rect 2010 2973 2013 3006
rect 2018 2996 2021 3023
rect 2026 3003 2029 3016
rect 2042 3013 2045 3073
rect 2074 3046 2077 3103
rect 2090 3053 2093 3116
rect 2098 3113 2117 3116
rect 2138 3113 2141 3143
rect 2098 3103 2101 3113
rect 2106 3103 2117 3106
rect 2074 3043 2085 3046
rect 2066 3013 2077 3016
rect 2082 3013 2085 3043
rect 2106 3013 2109 3086
rect 2114 3023 2133 3026
rect 2018 2993 2045 2996
rect 2018 2946 2021 2986
rect 1954 2853 2005 2856
rect 2010 2943 2021 2946
rect 1930 2813 1937 2816
rect 1954 2813 1957 2853
rect 2010 2836 2013 2943
rect 2002 2833 2013 2836
rect 1922 2773 1925 2806
rect 1934 2766 1937 2813
rect 1930 2763 1937 2766
rect 1914 2753 1921 2756
rect 1906 2703 1909 2726
rect 1918 2696 1921 2753
rect 1914 2693 1921 2696
rect 1842 2613 1845 2626
rect 1858 2613 1861 2626
rect 1834 2483 1837 2606
rect 1866 2576 1869 2606
rect 1882 2593 1885 2676
rect 1914 2626 1917 2693
rect 1914 2623 1921 2626
rect 1906 2576 1909 2616
rect 1866 2573 1909 2576
rect 1918 2566 1921 2623
rect 1930 2583 1933 2763
rect 1938 2713 1941 2736
rect 1946 2733 1949 2786
rect 1970 2743 1973 2806
rect 2002 2766 2005 2833
rect 2018 2813 2021 2936
rect 2026 2863 2029 2946
rect 2042 2923 2045 2993
rect 2050 2943 2053 3006
rect 2050 2826 2053 2936
rect 2058 2926 2061 3006
rect 2066 2966 2069 3006
rect 2074 2996 2077 3013
rect 2114 3003 2117 3023
rect 2122 2996 2125 3016
rect 2130 3013 2133 3023
rect 2074 2993 2125 2996
rect 2082 2973 2085 2986
rect 2122 2983 2125 2993
rect 2066 2963 2085 2966
rect 2066 2933 2069 2946
rect 2058 2923 2077 2926
rect 2082 2923 2085 2963
rect 2130 2943 2133 3006
rect 2138 2933 2141 3016
rect 2106 2923 2133 2926
rect 2074 2916 2077 2923
rect 2074 2913 2101 2916
rect 2122 2903 2125 2916
rect 2146 2886 2149 3136
rect 2170 3123 2173 3213
rect 2186 3133 2189 3196
rect 2154 3033 2157 3106
rect 2162 3026 2165 3066
rect 2154 3023 2165 3026
rect 2170 3023 2173 3056
rect 2194 3023 2197 3116
rect 2202 3113 2205 3196
rect 2218 3183 2221 3206
rect 2242 3176 2245 3216
rect 2298 3176 2301 3216
rect 2306 3203 2309 3216
rect 2314 3193 2317 3216
rect 2338 3183 2341 3226
rect 2386 3213 2389 3253
rect 2410 3176 2413 3253
rect 3074 3253 3117 3256
rect 2650 3233 2669 3236
rect 2674 3233 2685 3236
rect 2226 3173 2245 3176
rect 2258 3173 2301 3176
rect 2402 3173 2413 3176
rect 2226 3133 2229 3173
rect 2218 3113 2221 3126
rect 2226 3123 2237 3126
rect 2242 3083 2245 3136
rect 2258 3133 2261 3173
rect 2282 3143 2301 3146
rect 2282 3133 2285 3143
rect 2274 3113 2277 3126
rect 2226 3023 2253 3026
rect 2154 2933 2157 3023
rect 2178 3003 2181 3016
rect 2154 2916 2157 2926
rect 2162 2923 2165 2966
rect 2170 2916 2173 2936
rect 2154 2913 2173 2916
rect 2122 2883 2149 2886
rect 2050 2823 2061 2826
rect 2050 2766 2053 2816
rect 2058 2776 2061 2823
rect 2122 2813 2125 2883
rect 2178 2856 2181 2926
rect 2170 2853 2181 2856
rect 2170 2843 2173 2853
rect 2194 2846 2197 2936
rect 2202 2913 2205 3006
rect 2194 2843 2201 2846
rect 2074 2793 2077 2806
rect 2058 2773 2065 2776
rect 1978 2763 2005 2766
rect 2018 2763 2053 2766
rect 1962 2693 1965 2726
rect 1978 2603 1981 2763
rect 1986 2733 1989 2756
rect 2018 2723 2021 2763
rect 2034 2723 2037 2736
rect 2026 2646 2029 2706
rect 2062 2696 2065 2773
rect 2058 2693 2065 2696
rect 2026 2643 2037 2646
rect 2002 2616 2005 2626
rect 2034 2616 2037 2643
rect 2058 2623 2061 2693
rect 2074 2616 2077 2726
rect 2114 2723 2117 2806
rect 2154 2746 2157 2816
rect 2170 2793 2173 2806
rect 2198 2796 2201 2843
rect 2210 2813 2213 3016
rect 2226 2936 2229 3023
rect 2234 2946 2237 3016
rect 2266 3013 2269 3076
rect 2274 3013 2277 3106
rect 2282 3013 2293 3016
rect 2234 2943 2253 2946
rect 2226 2933 2237 2936
rect 2218 2913 2221 2926
rect 2226 2913 2229 2926
rect 2234 2903 2237 2933
rect 2242 2883 2245 2916
rect 2258 2906 2261 2936
rect 2266 2923 2269 3006
rect 2282 2993 2285 3006
rect 2290 2946 2293 3013
rect 2282 2943 2293 2946
rect 2282 2926 2285 2943
rect 2298 2926 2301 3136
rect 2306 3113 2309 3126
rect 2306 2983 2309 3036
rect 2314 3013 2317 3136
rect 2362 3133 2365 3146
rect 2322 3093 2325 3126
rect 2330 3106 2333 3126
rect 2330 3103 2341 3106
rect 2338 3056 2341 3103
rect 2330 3053 2341 3056
rect 2330 3033 2333 3053
rect 2274 2923 2285 2926
rect 2294 2923 2301 2926
rect 2258 2903 2277 2906
rect 2282 2893 2285 2916
rect 2294 2876 2297 2923
rect 2306 2886 2309 2946
rect 2322 2933 2325 2946
rect 2314 2903 2317 2916
rect 2306 2883 2317 2886
rect 2294 2873 2301 2876
rect 2194 2793 2201 2796
rect 2194 2776 2197 2793
rect 2170 2773 2197 2776
rect 2146 2743 2157 2746
rect 2122 2703 2125 2726
rect 2002 2613 2029 2616
rect 2034 2613 2061 2616
rect 2070 2613 2077 2616
rect 2002 2603 2013 2606
rect 1842 2563 1885 2566
rect 1918 2563 1925 2566
rect 1842 2533 1845 2563
rect 1858 2433 1861 2546
rect 1882 2523 1885 2563
rect 1810 2413 1817 2416
rect 1810 2393 1813 2413
rect 1730 2373 1749 2376
rect 1866 2373 1869 2466
rect 1922 2443 1925 2563
rect 1962 2533 1965 2546
rect 1930 2523 1941 2526
rect 2002 2523 2005 2603
rect 2010 2583 2013 2596
rect 2050 2586 2053 2606
rect 2050 2583 2061 2586
rect 2050 2536 2053 2583
rect 2070 2566 2073 2613
rect 2070 2563 2077 2566
rect 2074 2543 2077 2563
rect 2082 2546 2085 2606
rect 2114 2553 2117 2616
rect 2130 2613 2133 2626
rect 2082 2543 2109 2546
rect 2042 2533 2053 2536
rect 2082 2533 2085 2543
rect 2090 2533 2101 2536
rect 2106 2533 2109 2543
rect 2138 2536 2141 2736
rect 2146 2716 2149 2743
rect 2162 2736 2165 2746
rect 2154 2733 2165 2736
rect 2170 2716 2173 2773
rect 2250 2766 2253 2816
rect 2298 2813 2301 2873
rect 2314 2806 2317 2883
rect 2330 2856 2333 3026
rect 2338 3013 2357 3016
rect 2370 3013 2373 3036
rect 2378 3013 2381 3156
rect 2402 3133 2405 3173
rect 2434 3156 2437 3216
rect 2466 3193 2469 3206
rect 2474 3186 2477 3216
rect 2490 3203 2493 3226
rect 2514 3196 2517 3216
rect 2506 3193 2517 3196
rect 2474 3183 2493 3186
rect 2426 3153 2437 3156
rect 2410 3133 2413 3146
rect 2386 3103 2389 3126
rect 2402 3033 2405 3116
rect 2426 3103 2429 3153
rect 2418 3033 2421 3046
rect 2386 3013 2389 3026
rect 2434 3016 2437 3136
rect 2466 3133 2477 3136
rect 2482 3133 2485 3156
rect 2354 3006 2357 3013
rect 2338 2923 2341 3006
rect 2346 2983 2349 3006
rect 2354 3003 2365 3006
rect 2394 2996 2397 3016
rect 2402 3003 2405 3016
rect 2426 3013 2437 3016
rect 2362 2973 2365 2996
rect 2370 2993 2397 2996
rect 2346 2933 2349 2956
rect 2354 2893 2357 2966
rect 2370 2936 2373 2993
rect 2426 2956 2429 3013
rect 2442 2973 2445 3026
rect 2450 3013 2453 3026
rect 2466 3006 2469 3026
rect 2474 3013 2477 3126
rect 2482 3113 2485 3126
rect 2490 3093 2493 3183
rect 2506 3133 2509 3193
rect 2522 3123 2525 3136
rect 2530 3116 2533 3226
rect 2650 3223 2653 3233
rect 2666 3226 2669 3233
rect 2658 3216 2661 3226
rect 2666 3223 2685 3226
rect 2570 3193 2573 3216
rect 2466 3003 2477 3006
rect 2506 3003 2509 3116
rect 2514 3073 2517 3116
rect 2522 3113 2533 3116
rect 2538 3113 2541 3156
rect 2562 3123 2565 3166
rect 2594 3153 2597 3206
rect 2602 3143 2605 3216
rect 2610 3213 2621 3216
rect 2634 3213 2661 3216
rect 2618 3136 2621 3156
rect 2626 3146 2629 3206
rect 2650 3193 2653 3206
rect 2626 3143 2637 3146
rect 2570 3133 2589 3136
rect 2586 3113 2589 3133
rect 2602 3133 2613 3136
rect 2618 3133 2629 3136
rect 2522 3036 2525 3113
rect 2530 3103 2581 3106
rect 2518 3033 2525 3036
rect 2490 2993 2501 2996
rect 2426 2953 2453 2956
rect 2442 2936 2445 2946
rect 2362 2933 2373 2936
rect 2394 2933 2445 2936
rect 2362 2913 2365 2926
rect 2378 2863 2381 2926
rect 2394 2923 2397 2933
rect 2410 2923 2433 2926
rect 2442 2923 2445 2933
rect 2386 2903 2389 2916
rect 2394 2903 2397 2916
rect 2410 2913 2413 2923
rect 2418 2886 2421 2916
rect 2394 2883 2421 2886
rect 2430 2866 2433 2923
rect 2450 2916 2453 2953
rect 2442 2913 2453 2916
rect 2458 2913 2461 2926
rect 2466 2923 2469 2956
rect 2474 2933 2485 2936
rect 2490 2933 2493 2993
rect 2518 2976 2521 3033
rect 2530 3023 2565 3026
rect 2530 3003 2533 3023
rect 2538 3003 2541 3016
rect 2546 3013 2557 3016
rect 2562 3013 2565 3023
rect 2518 2973 2525 2976
rect 2546 2973 2549 3013
rect 2554 2993 2557 3006
rect 2562 2983 2565 3006
rect 2522 2933 2525 2973
rect 2570 2966 2573 3086
rect 2578 3003 2581 3103
rect 2602 3083 2605 3133
rect 2610 3113 2613 3126
rect 2586 3046 2589 3066
rect 2586 3043 2597 3046
rect 2594 2996 2597 3043
rect 2610 3023 2629 3026
rect 2610 3013 2613 3023
rect 2430 2863 2437 2866
rect 2330 2853 2341 2856
rect 2274 2793 2277 2806
rect 2306 2803 2317 2806
rect 2306 2776 2309 2803
rect 2306 2773 2333 2776
rect 2338 2773 2341 2853
rect 2234 2763 2253 2766
rect 2146 2713 2157 2716
rect 2154 2636 2157 2713
rect 2146 2633 2157 2636
rect 2166 2713 2173 2716
rect 2166 2636 2169 2713
rect 2166 2633 2173 2636
rect 2146 2613 2149 2633
rect 2146 2583 2149 2606
rect 2154 2593 2157 2616
rect 2170 2556 2173 2633
rect 2178 2603 2181 2736
rect 2194 2616 2197 2736
rect 2234 2706 2237 2763
rect 2226 2703 2237 2706
rect 2210 2666 2213 2686
rect 2186 2613 2197 2616
rect 2206 2663 2213 2666
rect 2114 2533 2141 2536
rect 2162 2553 2173 2556
rect 2042 2486 2045 2533
rect 2066 2513 2069 2526
rect 2042 2483 2053 2486
rect 2050 2463 2053 2483
rect 2058 2476 2061 2506
rect 2074 2493 2077 2526
rect 2090 2503 2093 2526
rect 2098 2523 2109 2526
rect 2114 2506 2117 2526
rect 2114 2503 2125 2506
rect 2058 2473 2069 2476
rect 1874 2423 1917 2426
rect 1874 2413 1877 2423
rect 1882 2403 1885 2416
rect 1890 2376 1893 2396
rect 1898 2383 1901 2416
rect 1914 2413 1917 2423
rect 1906 2376 1909 2406
rect 1890 2373 1909 2376
rect 1674 2333 1685 2336
rect 1714 2333 1733 2336
rect 1538 2243 1549 2246
rect 1490 2096 1493 2156
rect 1506 2153 1509 2196
rect 1514 2173 1517 2206
rect 1522 2193 1525 2216
rect 1530 2213 1533 2236
rect 1514 2133 1525 2136
rect 1490 2093 1501 2096
rect 1442 1793 1453 1796
rect 1410 1543 1413 1616
rect 1402 1523 1409 1526
rect 1406 1436 1409 1523
rect 1418 1513 1421 1646
rect 1426 1603 1429 1616
rect 1434 1586 1437 1736
rect 1442 1726 1445 1793
rect 1450 1733 1453 1766
rect 1442 1723 1453 1726
rect 1442 1603 1445 1676
rect 1434 1583 1441 1586
rect 1426 1496 1429 1556
rect 1438 1516 1441 1583
rect 1450 1533 1453 1723
rect 1458 1516 1461 1876
rect 1466 1773 1469 1826
rect 1466 1553 1469 1726
rect 1474 1553 1477 2006
rect 1482 1933 1485 2026
rect 1482 1636 1485 1916
rect 1490 1693 1493 2086
rect 1498 2033 1501 2093
rect 1506 2063 1509 2126
rect 1530 2123 1533 2166
rect 1538 2146 1541 2216
rect 1546 2156 1549 2243
rect 1546 2153 1557 2156
rect 1538 2143 1549 2146
rect 1530 2076 1533 2096
rect 1538 2083 1541 2136
rect 1546 2076 1549 2143
rect 1522 2073 1533 2076
rect 1538 2073 1549 2076
rect 1522 2026 1525 2073
rect 1522 2023 1533 2026
rect 1498 1943 1501 2006
rect 1514 1943 1517 2006
rect 1498 1863 1501 1936
rect 1506 1933 1517 1936
rect 1498 1793 1501 1836
rect 1506 1823 1509 1926
rect 1498 1663 1501 1736
rect 1506 1723 1509 1816
rect 1514 1813 1517 1926
rect 1522 1793 1525 1986
rect 1530 1923 1533 2023
rect 1538 2013 1541 2073
rect 1554 2043 1557 2153
rect 1562 2033 1565 2126
rect 1554 2016 1557 2026
rect 1554 2013 1565 2016
rect 1546 1983 1549 2006
rect 1554 1986 1557 2006
rect 1562 1996 1565 2013
rect 1570 2003 1573 2216
rect 1586 2146 1589 2226
rect 1578 2143 1589 2146
rect 1578 2003 1581 2143
rect 1594 2136 1597 2216
rect 1602 2156 1605 2226
rect 1610 2183 1613 2326
rect 1618 2163 1621 2196
rect 1602 2153 1621 2156
rect 1618 2143 1621 2153
rect 1626 2136 1629 2326
rect 1634 2323 1637 2333
rect 1642 2323 1653 2326
rect 1674 2323 1685 2326
rect 1634 2213 1637 2236
rect 1642 2213 1645 2266
rect 1650 2213 1653 2316
rect 1674 2306 1677 2323
rect 1666 2303 1677 2306
rect 1666 2236 1669 2303
rect 1666 2233 1677 2236
rect 1586 2133 1597 2136
rect 1562 1993 1573 1996
rect 1554 1983 1565 1986
rect 1554 1926 1557 1946
rect 1546 1923 1557 1926
rect 1530 1786 1533 1876
rect 1546 1846 1549 1923
rect 1562 1873 1565 1983
rect 1570 1933 1573 1993
rect 1546 1843 1557 1846
rect 1538 1803 1541 1826
rect 1522 1783 1533 1786
rect 1514 1733 1517 1746
rect 1522 1726 1525 1783
rect 1514 1723 1525 1726
rect 1514 1703 1517 1723
rect 1482 1633 1501 1636
rect 1482 1546 1485 1626
rect 1402 1433 1409 1436
rect 1422 1493 1429 1496
rect 1434 1513 1441 1516
rect 1450 1513 1461 1516
rect 1434 1493 1437 1513
rect 1402 1396 1405 1433
rect 1422 1426 1425 1493
rect 1422 1423 1429 1426
rect 1410 1403 1413 1416
rect 1426 1403 1429 1423
rect 1402 1393 1421 1396
rect 1402 1313 1405 1326
rect 1410 1323 1413 1386
rect 1418 1306 1421 1393
rect 1426 1313 1429 1336
rect 1414 1303 1421 1306
rect 1386 1123 1389 1296
rect 1394 1293 1405 1296
rect 1402 1226 1405 1293
rect 1398 1223 1405 1226
rect 1414 1226 1417 1303
rect 1434 1296 1437 1446
rect 1450 1336 1453 1513
rect 1466 1496 1469 1546
rect 1474 1543 1485 1546
rect 1462 1493 1469 1496
rect 1462 1356 1465 1493
rect 1462 1353 1469 1356
rect 1450 1333 1461 1336
rect 1442 1313 1453 1316
rect 1434 1293 1441 1296
rect 1414 1223 1421 1226
rect 1398 1146 1401 1223
rect 1394 1143 1401 1146
rect 1394 1016 1397 1143
rect 1402 1113 1405 1126
rect 1410 1043 1413 1206
rect 1394 1013 1405 1016
rect 1362 903 1365 916
rect 1370 863 1373 936
rect 1378 846 1381 946
rect 1374 843 1381 846
rect 1362 813 1365 826
rect 1374 776 1377 843
rect 1386 823 1389 956
rect 1394 913 1397 996
rect 1402 906 1405 1013
rect 1394 903 1405 906
rect 1386 803 1389 816
rect 1374 773 1381 776
rect 1378 753 1381 773
rect 1394 746 1397 903
rect 1410 863 1413 1006
rect 1402 803 1405 856
rect 1390 743 1397 746
rect 1362 723 1381 726
rect 1378 713 1381 723
rect 1390 686 1393 743
rect 1386 683 1393 686
rect 1402 683 1405 736
rect 1410 693 1413 816
rect 1362 563 1365 646
rect 1370 623 1373 666
rect 1370 543 1373 606
rect 1378 583 1381 606
rect 1386 526 1389 683
rect 1418 666 1421 1223
rect 1426 1213 1429 1276
rect 1426 1133 1429 1206
rect 1438 1146 1441 1293
rect 1434 1143 1441 1146
rect 1426 976 1429 1096
rect 1434 1003 1437 1143
rect 1450 1133 1453 1286
rect 1458 1176 1461 1333
rect 1466 1193 1469 1353
rect 1458 1173 1465 1176
rect 1462 1126 1465 1173
rect 1442 1013 1445 1126
rect 1458 1123 1465 1126
rect 1458 1056 1461 1123
rect 1458 1053 1465 1056
rect 1450 1023 1453 1046
rect 1426 973 1445 976
rect 1450 973 1453 1006
rect 1462 976 1465 1053
rect 1458 973 1465 976
rect 1426 893 1429 936
rect 1442 923 1445 973
rect 1450 906 1453 936
rect 1442 903 1453 906
rect 1426 706 1429 816
rect 1442 796 1445 903
rect 1442 793 1453 796
rect 1434 766 1437 776
rect 1450 766 1453 793
rect 1434 763 1453 766
rect 1434 723 1437 763
rect 1426 703 1437 706
rect 1410 663 1421 666
rect 1410 616 1413 663
rect 1434 626 1437 703
rect 1434 623 1445 626
rect 1450 623 1453 726
rect 1458 706 1461 973
rect 1474 956 1477 1536
rect 1482 1533 1493 1536
rect 1482 1423 1485 1466
rect 1490 1453 1493 1526
rect 1498 1506 1501 1633
rect 1506 1623 1509 1686
rect 1522 1586 1525 1606
rect 1518 1583 1525 1586
rect 1506 1533 1509 1546
rect 1518 1526 1521 1583
rect 1506 1513 1509 1526
rect 1518 1523 1525 1526
rect 1498 1503 1513 1506
rect 1482 1393 1485 1406
rect 1490 1393 1493 1446
rect 1482 1323 1485 1366
rect 1482 1283 1485 1316
rect 1482 1013 1485 1256
rect 1490 1196 1493 1316
rect 1498 1253 1501 1496
rect 1510 1436 1513 1503
rect 1522 1443 1525 1523
rect 1510 1433 1517 1436
rect 1506 1393 1509 1416
rect 1506 1333 1509 1366
rect 1498 1203 1501 1236
rect 1490 1193 1501 1196
rect 1490 1096 1493 1136
rect 1498 1113 1501 1193
rect 1490 1093 1497 1096
rect 1466 953 1477 956
rect 1466 896 1469 953
rect 1474 903 1477 946
rect 1466 893 1473 896
rect 1470 826 1473 893
rect 1470 823 1477 826
rect 1466 783 1469 806
rect 1466 723 1469 776
rect 1458 703 1465 706
rect 1378 523 1389 526
rect 1378 446 1381 523
rect 1378 443 1389 446
rect 1338 403 1357 406
rect 1338 333 1341 403
rect 1274 293 1277 316
rect 1306 313 1317 316
rect 1322 323 1333 326
rect 1262 233 1269 236
rect 1306 236 1309 313
rect 1322 246 1325 323
rect 1330 283 1333 316
rect 1354 313 1357 336
rect 1362 323 1365 426
rect 1370 273 1373 316
rect 1378 253 1381 406
rect 1386 266 1389 443
rect 1394 283 1397 616
rect 1410 613 1421 616
rect 1442 613 1445 623
rect 1462 616 1465 703
rect 1458 613 1465 616
rect 1410 516 1413 536
rect 1406 513 1413 516
rect 1406 436 1409 513
rect 1406 433 1413 436
rect 1402 323 1405 416
rect 1410 333 1413 433
rect 1418 413 1421 613
rect 1442 523 1445 606
rect 1426 493 1429 506
rect 1450 476 1453 556
rect 1458 513 1461 613
rect 1442 473 1453 476
rect 1442 426 1445 473
rect 1442 423 1453 426
rect 1450 403 1453 423
rect 1386 263 1397 266
rect 1322 243 1329 246
rect 1306 233 1317 236
rect 1250 193 1253 216
rect 1218 163 1229 166
rect 1262 166 1265 233
rect 1262 163 1269 166
rect 1218 146 1221 163
rect 1218 143 1261 146
rect 1258 133 1261 143
rect 1178 113 1205 116
rect 1250 33 1253 126
rect 1266 123 1269 163
rect 1274 133 1277 226
rect 1306 143 1309 216
rect 1314 193 1317 233
rect 1326 186 1329 243
rect 1346 243 1373 246
rect 1346 213 1349 243
rect 1354 213 1365 216
rect 1338 196 1341 206
rect 1346 203 1357 206
rect 1362 196 1365 206
rect 1338 193 1365 196
rect 1326 183 1349 186
rect 1346 133 1349 183
rect 1370 133 1373 243
rect 1378 193 1381 206
rect 1394 146 1397 263
rect 1386 143 1397 146
rect 1314 103 1317 126
rect 1338 83 1341 126
rect 1354 53 1357 126
rect 1386 123 1389 143
rect 1418 133 1421 326
rect 1426 313 1445 316
rect 1442 223 1445 313
rect 1458 293 1461 346
rect 1466 273 1469 526
rect 1474 523 1477 823
rect 1482 743 1485 996
rect 1494 986 1497 1093
rect 1506 1023 1509 1266
rect 1494 983 1509 986
rect 1490 933 1493 956
rect 1498 866 1501 976
rect 1490 863 1501 866
rect 1490 773 1493 863
rect 1498 813 1501 856
rect 1482 586 1485 656
rect 1490 603 1493 736
rect 1498 733 1501 806
rect 1506 626 1509 983
rect 1514 886 1517 1433
rect 1530 1423 1533 1726
rect 1538 1623 1541 1776
rect 1546 1733 1549 1756
rect 1546 1613 1549 1666
rect 1522 1383 1525 1406
rect 1530 1346 1533 1416
rect 1522 1343 1533 1346
rect 1522 1273 1525 1343
rect 1530 1293 1533 1336
rect 1522 1143 1525 1216
rect 1530 1183 1533 1226
rect 1530 1143 1533 1176
rect 1522 973 1525 1116
rect 1538 1063 1541 1606
rect 1554 1546 1557 1843
rect 1562 1823 1573 1826
rect 1578 1823 1581 1936
rect 1586 1923 1589 2133
rect 1594 2013 1597 2126
rect 1602 2093 1605 2136
rect 1610 2133 1629 2136
rect 1610 2086 1613 2133
rect 1606 2083 1613 2086
rect 1606 2026 1609 2083
rect 1602 2023 1609 2026
rect 1594 1923 1597 2006
rect 1602 1923 1605 2023
rect 1610 1993 1613 2006
rect 1618 1986 1621 2096
rect 1626 2033 1629 2106
rect 1610 1983 1621 1986
rect 1602 1896 1605 1916
rect 1594 1893 1605 1896
rect 1594 1836 1597 1893
rect 1594 1833 1605 1836
rect 1562 1573 1565 1646
rect 1554 1543 1565 1546
rect 1546 1533 1557 1536
rect 1546 1493 1549 1526
rect 1546 1333 1549 1406
rect 1554 1386 1557 1533
rect 1562 1403 1565 1543
rect 1570 1533 1573 1726
rect 1578 1603 1581 1796
rect 1586 1793 1589 1816
rect 1586 1686 1589 1746
rect 1586 1683 1597 1686
rect 1570 1506 1573 1526
rect 1578 1513 1581 1576
rect 1570 1503 1581 1506
rect 1570 1413 1573 1466
rect 1554 1383 1561 1386
rect 1578 1383 1581 1503
rect 1586 1423 1589 1683
rect 1602 1633 1605 1833
rect 1610 1813 1613 1983
rect 1618 1773 1621 1916
rect 1626 1816 1629 2016
rect 1634 2003 1637 2196
rect 1650 2096 1653 2166
rect 1658 2103 1661 2186
rect 1666 2113 1669 2216
rect 1650 2093 1669 2096
rect 1642 2003 1645 2076
rect 1650 1993 1653 2046
rect 1666 2013 1669 2093
rect 1658 2003 1669 2006
rect 1634 1903 1637 1936
rect 1642 1873 1645 1936
rect 1626 1813 1645 1816
rect 1626 1743 1629 1806
rect 1618 1676 1621 1736
rect 1634 1723 1637 1806
rect 1642 1803 1645 1813
rect 1650 1803 1653 1976
rect 1658 1943 1661 2003
rect 1610 1673 1621 1676
rect 1610 1633 1613 1673
rect 1594 1483 1597 1626
rect 1610 1616 1613 1626
rect 1602 1613 1613 1616
rect 1546 1303 1549 1326
rect 1546 1213 1549 1286
rect 1558 1246 1561 1383
rect 1586 1356 1589 1406
rect 1578 1353 1589 1356
rect 1570 1273 1573 1346
rect 1558 1243 1565 1246
rect 1546 1123 1549 1146
rect 1554 1106 1557 1236
rect 1550 1103 1557 1106
rect 1550 1036 1553 1103
rect 1550 1033 1557 1036
rect 1522 903 1525 946
rect 1530 923 1533 1016
rect 1546 993 1549 1006
rect 1554 936 1557 1033
rect 1562 1013 1565 1243
rect 1570 1123 1573 1206
rect 1570 996 1573 1026
rect 1546 933 1557 936
rect 1566 993 1573 996
rect 1566 926 1569 993
rect 1578 943 1581 1353
rect 1586 1313 1589 1346
rect 1594 1236 1597 1476
rect 1602 1323 1605 1586
rect 1610 1566 1613 1613
rect 1618 1583 1621 1636
rect 1626 1593 1629 1636
rect 1634 1573 1637 1636
rect 1610 1563 1617 1566
rect 1614 1506 1617 1563
rect 1626 1533 1629 1546
rect 1614 1503 1625 1506
rect 1610 1413 1613 1496
rect 1622 1446 1625 1503
rect 1622 1443 1629 1446
rect 1626 1423 1629 1443
rect 1618 1366 1621 1386
rect 1614 1363 1621 1366
rect 1614 1306 1617 1363
rect 1610 1303 1617 1306
rect 1594 1233 1601 1236
rect 1586 1173 1589 1226
rect 1598 1156 1601 1233
rect 1610 1206 1613 1303
rect 1626 1286 1629 1406
rect 1634 1403 1637 1526
rect 1622 1283 1629 1286
rect 1622 1226 1625 1283
rect 1634 1233 1637 1336
rect 1642 1313 1645 1766
rect 1658 1753 1661 1936
rect 1666 1773 1669 1956
rect 1674 1896 1677 2233
rect 1682 2043 1685 2316
rect 1722 2296 1725 2326
rect 1730 2303 1733 2333
rect 1746 2296 1749 2373
rect 1722 2293 1749 2296
rect 1770 2286 1773 2346
rect 1786 2293 1789 2346
rect 1834 2323 1837 2336
rect 1866 2323 1869 2366
rect 1874 2333 1877 2356
rect 1930 2343 1933 2406
rect 1922 2333 1933 2336
rect 1970 2326 1973 2386
rect 1978 2376 1981 2416
rect 2010 2403 2013 2416
rect 2034 2393 2037 2406
rect 2066 2396 2069 2473
rect 2058 2393 2069 2396
rect 1978 2373 2029 2376
rect 1986 2333 1989 2356
rect 2026 2333 2029 2373
rect 2034 2333 2037 2356
rect 1770 2283 1793 2286
rect 1706 2176 1709 2236
rect 1714 2206 1717 2276
rect 1722 2223 1733 2226
rect 1746 2213 1757 2216
rect 1714 2203 1725 2206
rect 1698 2136 1701 2176
rect 1706 2173 1717 2176
rect 1690 2133 1709 2136
rect 1698 2073 1701 2126
rect 1698 2003 1701 2056
rect 1682 1933 1685 1956
rect 1682 1916 1685 1926
rect 1690 1923 1693 1976
rect 1698 1923 1701 1946
rect 1706 1916 1709 2133
rect 1714 2096 1717 2173
rect 1722 2123 1725 2203
rect 1730 2193 1733 2206
rect 1730 2123 1733 2136
rect 1722 2113 1733 2116
rect 1714 2093 1725 2096
rect 1722 2026 1725 2093
rect 1738 2053 1741 2136
rect 1746 2103 1749 2213
rect 1714 2023 1725 2026
rect 1714 1953 1717 2023
rect 1722 1966 1725 2006
rect 1730 1973 1733 1996
rect 1722 1963 1733 1966
rect 1682 1913 1709 1916
rect 1674 1893 1681 1896
rect 1678 1836 1681 1893
rect 1674 1833 1681 1836
rect 1674 1756 1677 1833
rect 1690 1823 1693 1886
rect 1670 1753 1677 1756
rect 1650 1313 1653 1606
rect 1658 1503 1661 1746
rect 1670 1656 1673 1753
rect 1682 1743 1685 1816
rect 1698 1803 1701 1876
rect 1698 1776 1701 1796
rect 1694 1773 1701 1776
rect 1682 1703 1685 1726
rect 1694 1716 1697 1773
rect 1706 1723 1709 1806
rect 1694 1713 1701 1716
rect 1670 1653 1677 1656
rect 1674 1633 1677 1653
rect 1666 1583 1669 1606
rect 1674 1593 1677 1616
rect 1682 1603 1685 1686
rect 1690 1603 1693 1616
rect 1698 1596 1701 1713
rect 1714 1676 1717 1936
rect 1722 1923 1725 1936
rect 1730 1933 1733 1963
rect 1738 1916 1741 2006
rect 1746 1946 1749 2016
rect 1754 1956 1757 2206
rect 1762 2203 1765 2226
rect 1778 2213 1781 2236
rect 1790 2226 1793 2283
rect 1790 2223 1797 2226
rect 1762 2153 1789 2156
rect 1762 2143 1765 2153
rect 1762 2073 1765 2126
rect 1770 2103 1773 2136
rect 1778 2106 1781 2146
rect 1786 2133 1789 2153
rect 1778 2103 1789 2106
rect 1794 2056 1797 2223
rect 1802 2213 1805 2276
rect 1810 2223 1813 2246
rect 1778 2053 1797 2056
rect 1762 2003 1765 2016
rect 1770 2003 1773 2026
rect 1778 1986 1781 2053
rect 1770 1983 1781 1986
rect 1754 1953 1765 1956
rect 1746 1943 1757 1946
rect 1762 1943 1765 1953
rect 1730 1913 1741 1916
rect 1730 1846 1733 1913
rect 1746 1896 1749 1936
rect 1722 1843 1733 1846
rect 1742 1893 1749 1896
rect 1722 1733 1725 1843
rect 1742 1826 1745 1893
rect 1754 1873 1757 1943
rect 1762 1866 1765 1936
rect 1770 1933 1773 1983
rect 1778 1933 1781 1976
rect 1770 1903 1773 1926
rect 1778 1896 1781 1926
rect 1786 1916 1789 2046
rect 1794 2003 1797 2016
rect 1794 1973 1797 1996
rect 1794 1953 1797 1966
rect 1802 1946 1805 2206
rect 1826 2203 1829 2266
rect 1834 2146 1837 2316
rect 1874 2303 1877 2326
rect 1914 2306 1917 2326
rect 1970 2323 1989 2326
rect 1906 2303 1917 2306
rect 1906 2256 1909 2303
rect 1930 2296 1933 2316
rect 1970 2306 1973 2323
rect 1970 2303 1977 2306
rect 1930 2293 1941 2296
rect 1906 2253 1917 2256
rect 1842 2213 1845 2236
rect 1842 2153 1845 2206
rect 1858 2203 1861 2236
rect 1890 2233 1901 2236
rect 1874 2196 1877 2206
rect 1882 2203 1885 2216
rect 1898 2213 1901 2233
rect 1850 2193 1877 2196
rect 1794 1943 1805 1946
rect 1794 1923 1797 1943
rect 1810 1936 1813 2106
rect 1818 1973 1821 2146
rect 1834 2143 1869 2146
rect 1826 2133 1845 2136
rect 1826 2103 1829 2133
rect 1834 2096 1837 2126
rect 1826 2093 1837 2096
rect 1842 2123 1853 2126
rect 1802 1933 1813 1936
rect 1786 1913 1797 1916
rect 1778 1893 1785 1896
rect 1762 1863 1773 1866
rect 1738 1823 1745 1826
rect 1714 1673 1721 1676
rect 1706 1613 1709 1666
rect 1718 1626 1721 1673
rect 1714 1623 1721 1626
rect 1682 1593 1701 1596
rect 1658 1363 1661 1406
rect 1666 1343 1669 1516
rect 1658 1276 1661 1336
rect 1650 1273 1661 1276
rect 1666 1273 1669 1326
rect 1622 1223 1629 1226
rect 1610 1203 1621 1206
rect 1594 1153 1601 1156
rect 1514 883 1521 886
rect 1518 816 1521 883
rect 1514 813 1521 816
rect 1530 813 1533 826
rect 1546 813 1549 906
rect 1554 853 1557 926
rect 1566 923 1573 926
rect 1570 903 1573 923
rect 1514 766 1517 813
rect 1522 773 1525 796
rect 1514 763 1525 766
rect 1514 723 1517 736
rect 1522 643 1525 763
rect 1502 623 1509 626
rect 1482 583 1493 586
rect 1490 516 1493 583
rect 1502 526 1505 623
rect 1502 523 1509 526
rect 1482 513 1493 516
rect 1482 416 1485 513
rect 1506 503 1509 523
rect 1514 456 1517 616
rect 1506 453 1517 456
rect 1506 423 1509 453
rect 1522 433 1525 606
rect 1530 583 1533 706
rect 1538 653 1541 806
rect 1554 803 1557 816
rect 1570 783 1573 816
rect 1578 803 1581 916
rect 1546 743 1549 756
rect 1554 733 1557 746
rect 1562 723 1581 726
rect 1586 703 1589 1136
rect 1594 776 1597 1153
rect 1602 1076 1605 1136
rect 1610 1123 1613 1186
rect 1618 1096 1621 1203
rect 1626 1133 1629 1223
rect 1634 1133 1637 1216
rect 1650 1213 1653 1273
rect 1642 1203 1653 1206
rect 1666 1186 1669 1216
rect 1658 1183 1669 1186
rect 1658 1136 1661 1183
rect 1658 1133 1669 1136
rect 1626 1113 1629 1126
rect 1634 1106 1637 1126
rect 1634 1103 1645 1106
rect 1618 1093 1625 1096
rect 1602 1073 1613 1076
rect 1602 1013 1605 1066
rect 1610 1043 1613 1073
rect 1622 1036 1625 1093
rect 1642 1046 1645 1103
rect 1666 1096 1669 1133
rect 1618 1033 1625 1036
rect 1634 1043 1645 1046
rect 1658 1093 1669 1096
rect 1658 1046 1661 1093
rect 1658 1043 1669 1046
rect 1602 876 1605 976
rect 1610 893 1613 966
rect 1602 873 1609 876
rect 1606 816 1609 873
rect 1606 813 1613 816
rect 1602 793 1605 806
rect 1594 773 1601 776
rect 1530 513 1533 526
rect 1546 523 1549 606
rect 1554 503 1557 666
rect 1562 486 1565 656
rect 1558 483 1565 486
rect 1478 413 1485 416
rect 1478 366 1481 413
rect 1478 363 1485 366
rect 1474 323 1477 346
rect 1482 306 1485 363
rect 1490 336 1493 406
rect 1498 363 1501 406
rect 1506 363 1541 366
rect 1506 353 1509 363
rect 1522 343 1525 356
rect 1490 333 1501 336
rect 1478 303 1485 306
rect 1478 256 1481 303
rect 1498 286 1501 333
rect 1490 283 1501 286
rect 1490 263 1493 283
rect 1478 253 1485 256
rect 1482 226 1485 253
rect 1482 223 1489 226
rect 1498 223 1517 226
rect 1530 223 1533 336
rect 1538 323 1541 363
rect 1546 303 1549 416
rect 1558 356 1561 483
rect 1570 423 1573 696
rect 1578 433 1581 636
rect 1558 353 1565 356
rect 1570 353 1573 406
rect 1554 286 1557 336
rect 1562 306 1565 353
rect 1578 323 1581 396
rect 1562 303 1573 306
rect 1546 283 1557 286
rect 1546 236 1549 283
rect 1570 236 1573 303
rect 1546 233 1557 236
rect 1474 176 1477 216
rect 1466 173 1477 176
rect 1466 123 1469 173
rect 1486 166 1489 223
rect 1498 196 1501 206
rect 1514 203 1517 223
rect 1554 213 1557 233
rect 1562 233 1573 236
rect 1498 193 1525 196
rect 1482 163 1489 166
rect 1410 86 1413 116
rect 1482 113 1485 163
rect 1490 123 1493 136
rect 1538 113 1541 126
rect 1402 83 1413 86
rect 1546 83 1549 126
rect 1562 53 1565 233
rect 1578 183 1581 216
rect 1586 203 1589 676
rect 1598 656 1601 773
rect 1594 653 1601 656
rect 1594 623 1597 653
rect 1610 646 1613 813
rect 1618 796 1621 1033
rect 1626 973 1629 1006
rect 1626 933 1629 946
rect 1634 903 1637 1043
rect 1642 993 1645 1016
rect 1650 936 1653 1026
rect 1666 1016 1669 1043
rect 1642 933 1653 936
rect 1658 1013 1669 1016
rect 1642 876 1645 933
rect 1658 916 1661 1013
rect 1666 963 1669 1006
rect 1634 873 1645 876
rect 1654 913 1661 916
rect 1634 813 1637 873
rect 1654 826 1657 913
rect 1654 823 1661 826
rect 1666 823 1669 936
rect 1618 793 1629 796
rect 1626 726 1629 793
rect 1642 786 1645 816
rect 1618 723 1629 726
rect 1638 783 1645 786
rect 1618 703 1621 723
rect 1638 676 1641 783
rect 1650 723 1653 806
rect 1650 693 1653 716
rect 1638 673 1645 676
rect 1642 653 1645 673
rect 1610 643 1645 646
rect 1602 633 1629 636
rect 1602 546 1605 633
rect 1610 576 1613 626
rect 1626 613 1629 633
rect 1626 593 1629 606
rect 1610 573 1621 576
rect 1594 543 1605 546
rect 1594 493 1597 543
rect 1594 313 1597 426
rect 1602 346 1605 536
rect 1618 466 1621 573
rect 1634 563 1637 626
rect 1642 473 1645 643
rect 1610 463 1621 466
rect 1610 356 1613 463
rect 1626 423 1629 446
rect 1610 353 1629 356
rect 1602 343 1617 346
rect 1602 293 1605 336
rect 1614 276 1617 343
rect 1626 313 1629 353
rect 1634 306 1637 466
rect 1650 323 1653 626
rect 1658 606 1661 823
rect 1666 733 1669 816
rect 1666 673 1669 716
rect 1658 603 1669 606
rect 1666 536 1669 603
rect 1674 543 1677 1576
rect 1682 1433 1685 1593
rect 1682 1333 1685 1426
rect 1690 1333 1693 1556
rect 1698 1513 1701 1586
rect 1706 1493 1709 1526
rect 1706 1466 1709 1486
rect 1702 1463 1709 1466
rect 1714 1463 1717 1623
rect 1722 1593 1725 1606
rect 1722 1513 1725 1546
rect 1702 1366 1705 1463
rect 1714 1423 1717 1446
rect 1702 1363 1709 1366
rect 1682 1203 1685 1256
rect 1690 1196 1693 1246
rect 1682 1193 1693 1196
rect 1682 1003 1685 1193
rect 1698 1186 1701 1346
rect 1690 1183 1701 1186
rect 1690 1096 1693 1183
rect 1698 1116 1701 1166
rect 1706 1123 1709 1363
rect 1698 1113 1709 1116
rect 1690 1093 1701 1096
rect 1698 1036 1701 1093
rect 1690 1033 1701 1036
rect 1682 933 1685 946
rect 1682 783 1685 926
rect 1682 603 1685 756
rect 1682 536 1685 556
rect 1658 523 1661 536
rect 1666 533 1685 536
rect 1674 483 1677 516
rect 1682 466 1685 533
rect 1674 463 1685 466
rect 1674 406 1677 463
rect 1690 413 1693 1033
rect 1714 1016 1717 1406
rect 1722 1313 1725 1336
rect 1722 1273 1725 1306
rect 1722 1133 1725 1236
rect 1730 1196 1733 1816
rect 1738 1763 1741 1823
rect 1746 1813 1765 1816
rect 1746 1783 1749 1796
rect 1770 1793 1773 1863
rect 1782 1826 1785 1893
rect 1778 1823 1785 1826
rect 1778 1786 1781 1823
rect 1754 1783 1781 1786
rect 1738 1593 1741 1656
rect 1738 1543 1741 1586
rect 1738 1523 1741 1536
rect 1746 1443 1749 1626
rect 1738 1326 1741 1336
rect 1746 1333 1749 1346
rect 1754 1336 1757 1783
rect 1786 1776 1789 1806
rect 1762 1773 1789 1776
rect 1762 1713 1765 1773
rect 1770 1616 1773 1746
rect 1762 1613 1773 1616
rect 1778 1613 1781 1636
rect 1762 1346 1765 1613
rect 1770 1586 1773 1606
rect 1770 1583 1777 1586
rect 1774 1426 1777 1583
rect 1786 1533 1789 1716
rect 1794 1603 1797 1913
rect 1802 1883 1805 1933
rect 1818 1926 1821 1956
rect 1826 1946 1829 2093
rect 1842 2086 1845 2123
rect 1858 2113 1861 2136
rect 1834 2083 1845 2086
rect 1834 2063 1837 2083
rect 1850 2073 1861 2076
rect 1850 2023 1853 2073
rect 1834 1953 1837 1976
rect 1842 1963 1845 2006
rect 1858 1946 1861 2036
rect 1866 2026 1869 2143
rect 1874 2116 1877 2186
rect 1882 2133 1885 2146
rect 1890 2126 1893 2206
rect 1898 2153 1901 2206
rect 1882 2123 1901 2126
rect 1874 2113 1893 2116
rect 1874 2033 1877 2106
rect 1866 2023 1877 2026
rect 1826 1943 1845 1946
rect 1810 1923 1821 1926
rect 1810 1876 1813 1916
rect 1826 1906 1829 1936
rect 1834 1923 1837 1936
rect 1806 1873 1813 1876
rect 1822 1903 1829 1906
rect 1806 1766 1809 1873
rect 1822 1846 1825 1903
rect 1822 1843 1829 1846
rect 1818 1813 1821 1826
rect 1802 1763 1809 1766
rect 1802 1716 1805 1763
rect 1810 1723 1813 1746
rect 1818 1733 1821 1806
rect 1802 1713 1813 1716
rect 1802 1623 1805 1646
rect 1802 1586 1805 1606
rect 1794 1583 1805 1586
rect 1794 1533 1797 1583
rect 1810 1553 1813 1713
rect 1770 1423 1777 1426
rect 1770 1363 1773 1423
rect 1786 1413 1789 1526
rect 1762 1343 1773 1346
rect 1754 1333 1765 1336
rect 1738 1323 1757 1326
rect 1762 1306 1765 1333
rect 1758 1303 1765 1306
rect 1738 1223 1741 1236
rect 1746 1233 1749 1256
rect 1738 1213 1749 1216
rect 1758 1206 1761 1303
rect 1770 1213 1773 1343
rect 1754 1203 1761 1206
rect 1730 1193 1741 1196
rect 1722 1083 1725 1126
rect 1738 1086 1741 1193
rect 1754 1186 1757 1203
rect 1730 1083 1741 1086
rect 1750 1183 1757 1186
rect 1762 1193 1773 1196
rect 1750 1086 1753 1183
rect 1750 1083 1757 1086
rect 1706 1013 1717 1016
rect 1706 933 1709 1013
rect 1714 986 1717 1006
rect 1714 983 1721 986
rect 1698 733 1701 926
rect 1706 903 1709 916
rect 1706 823 1709 896
rect 1718 886 1721 983
rect 1714 883 1721 886
rect 1698 523 1701 536
rect 1698 423 1701 446
rect 1706 423 1709 776
rect 1714 623 1717 883
rect 1722 803 1725 866
rect 1722 783 1725 796
rect 1722 723 1725 776
rect 1730 656 1733 1083
rect 1746 1023 1749 1066
rect 1738 913 1741 1016
rect 1746 973 1749 1016
rect 1738 813 1741 826
rect 1746 796 1749 926
rect 1742 793 1749 796
rect 1742 706 1745 793
rect 1738 703 1745 706
rect 1738 683 1741 703
rect 1730 653 1737 656
rect 1722 613 1725 646
rect 1734 606 1737 653
rect 1730 603 1737 606
rect 1746 603 1749 696
rect 1754 656 1757 1083
rect 1762 753 1765 1193
rect 1778 1153 1781 1406
rect 1786 1223 1789 1326
rect 1794 1293 1797 1366
rect 1770 1143 1781 1146
rect 1786 1056 1789 1216
rect 1794 1123 1797 1256
rect 1770 853 1773 1056
rect 1786 1053 1797 1056
rect 1794 1013 1797 1053
rect 1778 1003 1797 1006
rect 1794 993 1797 1003
rect 1778 906 1781 986
rect 1786 983 1797 986
rect 1786 923 1789 983
rect 1778 903 1785 906
rect 1794 903 1797 936
rect 1802 933 1805 1536
rect 1818 1523 1821 1606
rect 1826 1506 1829 1843
rect 1834 1763 1837 1916
rect 1842 1913 1845 1943
rect 1850 1943 1861 1946
rect 1842 1826 1845 1906
rect 1850 1836 1853 1943
rect 1866 1936 1869 2016
rect 1874 2003 1877 2023
rect 1858 1926 1861 1936
rect 1866 1933 1877 1936
rect 1882 1933 1885 1956
rect 1858 1923 1869 1926
rect 1858 1843 1861 1916
rect 1866 1873 1869 1923
rect 1874 1913 1877 1933
rect 1890 1926 1893 2113
rect 1906 2023 1909 2226
rect 1914 1996 1917 2253
rect 1938 2246 1941 2293
rect 1930 2243 1941 2246
rect 1930 2206 1933 2243
rect 1954 2213 1957 2226
rect 1922 2203 1933 2206
rect 1922 2116 1925 2203
rect 1930 2173 1933 2196
rect 1962 2193 1965 2286
rect 1974 2226 1977 2303
rect 1970 2223 1977 2226
rect 1946 2136 1949 2156
rect 1954 2143 1965 2146
rect 1938 2133 1957 2136
rect 1922 2113 1933 2116
rect 1930 2066 1933 2113
rect 1954 2073 1957 2126
rect 1922 2063 1933 2066
rect 1922 2043 1925 2063
rect 1922 2033 1957 2036
rect 1922 2003 1925 2033
rect 1946 2016 1949 2026
rect 1930 2013 1949 2016
rect 1914 1993 1925 1996
rect 1898 1933 1901 1976
rect 1906 1933 1917 1936
rect 1890 1923 1901 1926
rect 1906 1923 1917 1926
rect 1882 1876 1885 1896
rect 1878 1873 1885 1876
rect 1850 1833 1861 1836
rect 1842 1823 1853 1826
rect 1850 1813 1853 1823
rect 1842 1803 1853 1806
rect 1858 1803 1861 1833
rect 1866 1803 1869 1826
rect 1850 1733 1853 1803
rect 1878 1796 1881 1873
rect 1878 1793 1885 1796
rect 1882 1776 1885 1793
rect 1866 1773 1885 1776
rect 1866 1723 1869 1773
rect 1834 1696 1837 1716
rect 1834 1693 1845 1696
rect 1842 1636 1845 1693
rect 1834 1633 1845 1636
rect 1834 1603 1837 1633
rect 1822 1503 1829 1506
rect 1834 1503 1837 1536
rect 1842 1533 1845 1616
rect 1850 1533 1853 1566
rect 1858 1553 1861 1656
rect 1866 1613 1869 1686
rect 1874 1566 1877 1766
rect 1882 1666 1885 1773
rect 1890 1673 1893 1923
rect 1906 1913 1909 1923
rect 1898 1826 1901 1846
rect 1898 1823 1905 1826
rect 1902 1756 1905 1823
rect 1898 1753 1905 1756
rect 1898 1733 1901 1753
rect 1882 1663 1893 1666
rect 1890 1653 1893 1663
rect 1898 1653 1901 1726
rect 1914 1723 1917 1906
rect 1922 1813 1925 1993
rect 1930 1893 1933 2013
rect 1938 1943 1941 2006
rect 1938 1886 1941 1936
rect 1930 1883 1941 1886
rect 1930 1743 1933 1883
rect 1938 1823 1941 1846
rect 1938 1736 1941 1806
rect 1930 1733 1941 1736
rect 1930 1716 1933 1733
rect 1930 1713 1941 1716
rect 1938 1696 1941 1713
rect 1934 1693 1941 1696
rect 1906 1646 1909 1686
rect 1882 1643 1909 1646
rect 1882 1603 1885 1643
rect 1874 1563 1885 1566
rect 1842 1523 1853 1526
rect 1858 1523 1861 1546
rect 1810 1413 1813 1436
rect 1810 1133 1813 1336
rect 1822 1276 1825 1503
rect 1822 1273 1829 1276
rect 1826 1253 1829 1273
rect 1834 1246 1837 1496
rect 1850 1423 1853 1523
rect 1866 1493 1869 1556
rect 1850 1383 1853 1406
rect 1858 1393 1861 1406
rect 1866 1366 1869 1456
rect 1858 1363 1869 1366
rect 1874 1363 1877 1556
rect 1850 1326 1853 1346
rect 1818 1243 1837 1246
rect 1846 1323 1853 1326
rect 1846 1246 1849 1323
rect 1846 1243 1853 1246
rect 1818 1223 1821 1243
rect 1818 1146 1821 1216
rect 1826 1166 1829 1243
rect 1834 1176 1837 1236
rect 1850 1213 1853 1243
rect 1850 1176 1853 1186
rect 1834 1173 1853 1176
rect 1858 1173 1861 1363
rect 1882 1356 1885 1563
rect 1890 1553 1893 1636
rect 1898 1613 1901 1636
rect 1934 1626 1937 1693
rect 1906 1623 1917 1626
rect 1906 1613 1909 1623
rect 1898 1546 1901 1556
rect 1914 1546 1917 1623
rect 1922 1553 1925 1626
rect 1930 1623 1937 1626
rect 1890 1543 1901 1546
rect 1890 1403 1893 1543
rect 1898 1523 1901 1536
rect 1906 1533 1909 1546
rect 1914 1543 1925 1546
rect 1922 1526 1925 1543
rect 1930 1533 1933 1623
rect 1906 1506 1909 1526
rect 1914 1516 1917 1526
rect 1922 1523 1933 1526
rect 1938 1523 1941 1616
rect 1914 1513 1941 1516
rect 1906 1503 1933 1506
rect 1866 1353 1885 1356
rect 1866 1256 1869 1353
rect 1874 1343 1885 1346
rect 1874 1273 1877 1326
rect 1890 1273 1893 1336
rect 1898 1323 1901 1446
rect 1906 1313 1909 1406
rect 1866 1253 1873 1256
rect 1826 1163 1837 1166
rect 1818 1143 1825 1146
rect 1822 1086 1825 1143
rect 1834 1096 1837 1163
rect 1850 1103 1853 1173
rect 1870 1136 1873 1253
rect 1870 1133 1877 1136
rect 1834 1093 1853 1096
rect 1822 1083 1845 1086
rect 1810 1056 1813 1076
rect 1810 1053 1821 1056
rect 1818 986 1821 1053
rect 1810 983 1821 986
rect 1810 916 1813 983
rect 1834 973 1837 1026
rect 1842 1016 1845 1083
rect 1850 1033 1853 1093
rect 1842 1013 1849 1016
rect 1818 933 1821 966
rect 1834 933 1837 966
rect 1846 926 1849 1013
rect 1858 963 1861 1026
rect 1866 1013 1869 1126
rect 1866 946 1869 1006
rect 1806 913 1813 916
rect 1762 673 1765 736
rect 1770 723 1773 806
rect 1782 796 1785 903
rect 1806 836 1809 913
rect 1818 843 1821 926
rect 1826 913 1829 926
rect 1842 923 1849 926
rect 1858 943 1869 946
rect 1806 833 1813 836
rect 1794 803 1797 816
rect 1778 793 1785 796
rect 1778 706 1781 793
rect 1786 743 1789 776
rect 1802 773 1805 816
rect 1802 716 1805 736
rect 1810 733 1813 833
rect 1842 826 1845 923
rect 1858 836 1861 943
rect 1874 853 1877 1133
rect 1882 906 1885 1256
rect 1890 1113 1893 1226
rect 1906 1223 1909 1236
rect 1906 1176 1909 1216
rect 1914 1206 1917 1496
rect 1922 1376 1925 1426
rect 1930 1406 1933 1503
rect 1946 1463 1949 2006
rect 1954 2003 1957 2033
rect 1954 1953 1957 1996
rect 1962 1983 1965 2126
rect 1970 2086 1973 2223
rect 1978 2193 1981 2206
rect 1978 2123 1981 2176
rect 1970 2083 1981 2086
rect 1954 1916 1957 1936
rect 1970 1923 1973 2076
rect 1978 1946 1981 2083
rect 1986 2073 1989 2276
rect 1994 2133 1997 2296
rect 2002 2223 2005 2266
rect 2026 2246 2029 2326
rect 2058 2323 2061 2393
rect 2082 2376 2085 2416
rect 2114 2413 2117 2496
rect 2122 2423 2125 2503
rect 2130 2483 2133 2526
rect 2146 2513 2149 2526
rect 2162 2506 2165 2553
rect 2186 2533 2189 2613
rect 2206 2606 2209 2663
rect 2226 2646 2229 2703
rect 2242 2686 2245 2726
rect 2274 2723 2277 2766
rect 2282 2733 2285 2746
rect 2242 2683 2277 2686
rect 2218 2643 2229 2646
rect 2218 2613 2221 2643
rect 2274 2626 2277 2683
rect 2306 2653 2309 2726
rect 2330 2703 2333 2773
rect 2338 2733 2341 2756
rect 2346 2713 2349 2736
rect 2354 2723 2357 2816
rect 2418 2813 2421 2836
rect 2434 2826 2437 2863
rect 2442 2833 2445 2913
rect 2482 2906 2485 2926
rect 2450 2903 2485 2906
rect 2506 2903 2509 2926
rect 2546 2913 2549 2926
rect 2554 2886 2557 2966
rect 2546 2883 2557 2886
rect 2566 2963 2573 2966
rect 2590 2993 2597 2996
rect 2434 2823 2461 2826
rect 2370 2793 2373 2806
rect 2362 2723 2373 2726
rect 2266 2623 2277 2626
rect 2206 2603 2213 2606
rect 2234 2603 2237 2616
rect 2210 2586 2213 2603
rect 2210 2583 2229 2586
rect 2226 2536 2229 2583
rect 2266 2576 2269 2623
rect 2266 2573 2277 2576
rect 2218 2533 2229 2536
rect 2162 2503 2173 2506
rect 2162 2456 2165 2486
rect 2170 2473 2173 2503
rect 2162 2453 2169 2456
rect 2138 2393 2141 2436
rect 2082 2373 2093 2376
rect 2090 2333 2093 2373
rect 2106 2333 2125 2336
rect 2154 2333 2157 2396
rect 2166 2346 2169 2453
rect 2218 2446 2221 2533
rect 2218 2443 2229 2446
rect 2162 2343 2169 2346
rect 2018 2243 2029 2246
rect 2002 2136 2005 2216
rect 2010 2143 2013 2166
rect 2002 2133 2013 2136
rect 1986 2006 1989 2046
rect 2002 2036 2005 2133
rect 2018 2116 2021 2243
rect 2026 2183 2029 2236
rect 1994 2033 2005 2036
rect 2014 2113 2021 2116
rect 2014 2036 2017 2113
rect 2014 2033 2021 2036
rect 1994 2013 1997 2033
rect 2002 2013 2013 2016
rect 1986 2003 2005 2006
rect 1978 1943 1989 1946
rect 1954 1913 1961 1916
rect 1958 1846 1961 1913
rect 1978 1906 1981 1936
rect 1986 1933 1989 1943
rect 1994 1933 1997 1966
rect 1954 1843 1961 1846
rect 1974 1903 1981 1906
rect 1954 1753 1957 1843
rect 1974 1826 1977 1903
rect 1962 1803 1965 1826
rect 1974 1823 1981 1826
rect 1978 1806 1981 1823
rect 1970 1803 1981 1806
rect 1986 1803 1989 1926
rect 1994 1883 1997 1926
rect 1954 1613 1957 1746
rect 1962 1716 1965 1736
rect 1970 1733 1973 1803
rect 1986 1736 1989 1786
rect 1982 1733 1989 1736
rect 1962 1713 1973 1716
rect 1970 1636 1973 1713
rect 1962 1633 1973 1636
rect 1962 1613 1965 1633
rect 1982 1626 1985 1733
rect 1994 1626 1997 1726
rect 2002 1703 2005 2003
rect 2010 1963 2013 2006
rect 2018 1973 2021 2033
rect 2018 1926 2021 1936
rect 2026 1933 2029 2136
rect 2034 2103 2037 2256
rect 2042 2223 2045 2246
rect 2042 2143 2045 2206
rect 2042 2093 2045 2126
rect 2050 2106 2053 2316
rect 2090 2253 2093 2316
rect 2098 2236 2101 2326
rect 2058 2233 2101 2236
rect 2058 2193 2061 2233
rect 2058 2123 2061 2166
rect 2066 2133 2069 2216
rect 2074 2193 2077 2216
rect 2098 2213 2101 2233
rect 2098 2196 2101 2206
rect 2082 2193 2101 2196
rect 2082 2123 2085 2136
rect 2098 2126 2101 2176
rect 2090 2123 2101 2126
rect 2050 2103 2057 2106
rect 2034 2023 2037 2066
rect 2010 1923 2021 1926
rect 2034 1923 2037 2006
rect 2010 1893 2013 1923
rect 2042 1916 2045 2076
rect 2054 2036 2057 2103
rect 2066 2083 2069 2116
rect 2050 2033 2057 2036
rect 2050 1986 2053 2033
rect 2058 2003 2061 2016
rect 2074 2013 2077 2036
rect 2050 1983 2069 1986
rect 2018 1913 2045 1916
rect 2018 1813 2021 1906
rect 2050 1826 2053 1936
rect 2058 1903 2061 1976
rect 2034 1783 2037 1826
rect 2046 1823 2053 1826
rect 2046 1756 2049 1823
rect 2034 1753 2049 1756
rect 2010 1723 2013 1746
rect 2018 1723 2021 1736
rect 2010 1626 2013 1636
rect 1982 1623 1989 1626
rect 1994 1623 2013 1626
rect 1954 1593 1957 1606
rect 1978 1596 1981 1606
rect 1962 1593 1981 1596
rect 1954 1533 1957 1546
rect 1962 1526 1965 1593
rect 1954 1523 1965 1526
rect 1954 1473 1957 1523
rect 1946 1423 1949 1456
rect 1962 1423 1965 1516
rect 1970 1453 1973 1566
rect 1978 1523 1981 1586
rect 1986 1446 1989 1623
rect 1994 1533 1997 1616
rect 2002 1563 2005 1616
rect 2010 1583 2013 1616
rect 2026 1603 2029 1686
rect 2034 1603 2037 1753
rect 2058 1746 2061 1816
rect 2066 1803 2069 1983
rect 2042 1733 2045 1746
rect 2050 1743 2061 1746
rect 2050 1723 2053 1736
rect 2002 1446 2005 1536
rect 2010 1503 2013 1526
rect 2018 1506 2021 1536
rect 2026 1533 2029 1586
rect 2034 1533 2037 1546
rect 2026 1513 2029 1526
rect 2018 1503 2029 1506
rect 1986 1443 1997 1446
rect 2002 1443 2021 1446
rect 1954 1413 1973 1416
rect 1930 1403 1949 1406
rect 1962 1386 1965 1406
rect 1970 1393 1973 1413
rect 1978 1403 1981 1416
rect 1962 1383 1981 1386
rect 1922 1373 1965 1376
rect 1938 1343 1957 1346
rect 1938 1333 1941 1343
rect 1922 1303 1925 1326
rect 1922 1223 1925 1276
rect 1914 1203 1921 1206
rect 1898 1173 1909 1176
rect 1898 1113 1901 1173
rect 1906 1106 1909 1156
rect 1898 1103 1909 1106
rect 1898 1026 1901 1103
rect 1918 1096 1921 1203
rect 1890 1023 1901 1026
rect 1914 1093 1921 1096
rect 1890 943 1893 1023
rect 1898 1003 1909 1006
rect 1914 986 1917 1093
rect 1906 983 1917 986
rect 1890 923 1893 936
rect 1882 903 1893 906
rect 1858 833 1869 836
rect 1834 823 1845 826
rect 1818 783 1821 806
rect 1818 726 1821 776
rect 1798 713 1805 716
rect 1810 723 1821 726
rect 1774 703 1781 706
rect 1754 653 1761 656
rect 1730 533 1733 603
rect 1758 596 1761 653
rect 1774 636 1777 703
rect 1774 633 1781 636
rect 1770 603 1773 616
rect 1754 593 1761 596
rect 1714 456 1717 526
rect 1730 473 1733 526
rect 1738 456 1741 536
rect 1714 453 1741 456
rect 1738 413 1741 426
rect 1746 413 1749 516
rect 1754 406 1757 593
rect 1778 526 1781 633
rect 1786 603 1789 706
rect 1798 646 1801 713
rect 1798 643 1805 646
rect 1794 593 1797 626
rect 1774 523 1781 526
rect 1762 423 1765 486
rect 1774 426 1777 523
rect 1774 423 1781 426
rect 1674 403 1685 406
rect 1658 333 1661 356
rect 1610 273 1617 276
rect 1630 303 1637 306
rect 1594 183 1597 256
rect 1570 113 1581 116
rect 1610 96 1613 273
rect 1630 246 1633 303
rect 1642 253 1645 316
rect 1626 243 1633 246
rect 1626 223 1629 243
rect 1666 233 1669 326
rect 1674 323 1677 336
rect 1682 323 1685 403
rect 1650 223 1661 226
rect 1626 213 1653 216
rect 1626 103 1629 213
rect 1658 173 1661 223
rect 1634 96 1637 116
rect 1610 93 1637 96
rect 1642 86 1645 126
rect 1666 103 1669 226
rect 1674 173 1677 296
rect 1714 246 1717 266
rect 1706 243 1717 246
rect 1706 196 1709 243
rect 1730 233 1733 336
rect 1738 306 1741 406
rect 1746 403 1757 406
rect 1778 403 1781 423
rect 1786 403 1789 516
rect 1802 506 1805 643
rect 1810 603 1813 723
rect 1834 716 1837 823
rect 1850 813 1861 816
rect 1850 776 1853 813
rect 1858 796 1861 806
rect 1866 803 1869 833
rect 1890 826 1893 903
rect 1906 896 1909 983
rect 1922 923 1925 1006
rect 1930 1003 1933 1326
rect 1954 1303 1957 1343
rect 1962 1286 1965 1373
rect 1954 1283 1965 1286
rect 1938 1196 1941 1266
rect 1938 1193 1945 1196
rect 1942 1136 1945 1193
rect 1954 1146 1957 1283
rect 1970 1206 1973 1366
rect 1978 1213 1981 1383
rect 1962 1183 1965 1206
rect 1970 1203 1977 1206
rect 1954 1143 1965 1146
rect 1942 1133 1957 1136
rect 1938 936 1941 1126
rect 1946 1013 1949 1026
rect 1930 933 1941 936
rect 1938 903 1941 926
rect 1946 923 1949 986
rect 1906 893 1941 896
rect 1938 836 1941 893
rect 1954 836 1957 1133
rect 1962 1123 1965 1143
rect 1974 1096 1977 1203
rect 1986 1103 1989 1443
rect 1994 1213 1997 1416
rect 2002 1333 2005 1436
rect 2010 1413 2013 1426
rect 2018 1413 2021 1443
rect 2010 1403 2021 1406
rect 2010 1323 2013 1386
rect 2026 1376 2029 1503
rect 2034 1433 2037 1526
rect 2042 1513 2045 1716
rect 2050 1623 2053 1646
rect 2058 1613 2061 1706
rect 2034 1403 2037 1426
rect 2042 1413 2045 1446
rect 2018 1373 2029 1376
rect 2018 1316 2021 1373
rect 2034 1333 2037 1396
rect 2010 1313 2021 1316
rect 1994 1113 1997 1136
rect 2002 1103 2005 1256
rect 1974 1093 1981 1096
rect 1962 933 1965 996
rect 1978 976 1981 1093
rect 2002 1003 2005 1026
rect 2010 1013 2013 1313
rect 2018 1236 2021 1296
rect 2026 1253 2029 1316
rect 2018 1233 2025 1236
rect 2034 1233 2037 1326
rect 2042 1323 2045 1386
rect 2022 1146 2025 1233
rect 2018 1143 2025 1146
rect 1974 973 1981 976
rect 1974 906 1977 973
rect 1986 913 1989 966
rect 1974 903 1981 906
rect 1938 833 1949 836
rect 1954 833 1973 836
rect 1890 823 1909 826
rect 1874 796 1877 816
rect 1858 793 1877 796
rect 1850 773 1861 776
rect 1850 723 1853 746
rect 1834 713 1845 716
rect 1818 523 1821 646
rect 1834 613 1837 646
rect 1842 613 1845 713
rect 1842 546 1845 606
rect 1842 543 1853 546
rect 1842 523 1845 536
rect 1802 503 1813 506
rect 1810 416 1813 503
rect 1842 443 1845 516
rect 1850 513 1853 543
rect 1802 413 1813 416
rect 1746 323 1749 403
rect 1762 313 1765 386
rect 1738 303 1749 306
rect 1746 246 1749 303
rect 1794 296 1797 326
rect 1778 293 1797 296
rect 1746 243 1757 246
rect 1730 203 1733 216
rect 1754 213 1757 243
rect 1706 193 1717 196
rect 1690 133 1693 176
rect 1714 143 1717 193
rect 1738 133 1741 206
rect 1754 146 1757 206
rect 1778 166 1781 293
rect 1802 276 1805 413
rect 1810 393 1837 396
rect 1834 386 1837 393
rect 1834 383 1845 386
rect 1818 323 1821 346
rect 1834 323 1837 383
rect 1850 316 1853 406
rect 1858 396 1861 773
rect 1874 633 1877 726
rect 1866 603 1869 616
rect 1874 603 1877 626
rect 1890 616 1893 816
rect 1906 766 1909 823
rect 1930 783 1933 806
rect 1898 743 1901 766
rect 1906 763 1917 766
rect 1914 646 1917 763
rect 1938 733 1941 816
rect 1938 693 1941 726
rect 1906 643 1917 646
rect 1906 626 1909 643
rect 1882 613 1893 616
rect 1902 623 1909 626
rect 1866 503 1869 526
rect 1882 426 1885 613
rect 1890 563 1893 606
rect 1902 536 1905 623
rect 1930 616 1933 626
rect 1930 613 1941 616
rect 1914 603 1925 606
rect 1946 603 1949 833
rect 1962 816 1965 826
rect 1954 813 1965 816
rect 1970 756 1973 833
rect 1954 753 1973 756
rect 1954 703 1957 753
rect 1962 723 1965 746
rect 1902 533 1909 536
rect 1914 533 1917 603
rect 1954 596 1957 636
rect 1970 626 1973 736
rect 1978 723 1981 903
rect 1994 863 1997 946
rect 2002 933 2005 996
rect 2018 923 2021 1143
rect 2034 1133 2037 1186
rect 2026 1063 2029 1126
rect 2026 1013 2029 1026
rect 2026 963 2029 1006
rect 2034 1003 2037 1116
rect 2026 903 2029 936
rect 2034 886 2037 926
rect 2026 883 2037 886
rect 1986 803 1989 856
rect 2026 826 2029 883
rect 2042 853 2045 1316
rect 2050 946 2053 1606
rect 2066 1603 2069 1726
rect 2058 1526 2061 1586
rect 2066 1533 2069 1596
rect 2058 1523 2069 1526
rect 2074 1523 2077 1976
rect 2082 1943 2085 2116
rect 2090 2093 2093 2123
rect 2106 2116 2109 2206
rect 2114 2203 2117 2286
rect 2122 2213 2125 2333
rect 2122 2193 2125 2206
rect 2098 2113 2109 2116
rect 2098 2073 2101 2113
rect 2106 2076 2109 2106
rect 2114 2083 2117 2116
rect 2122 2076 2125 2186
rect 2130 2173 2133 2246
rect 2138 2203 2141 2216
rect 2146 2203 2149 2236
rect 2106 2073 2125 2076
rect 2090 1983 2093 2016
rect 2098 1966 2101 2036
rect 2114 2006 2117 2016
rect 2106 2003 2117 2006
rect 2106 1973 2109 2003
rect 2114 1966 2117 1996
rect 2122 1993 2125 2016
rect 2098 1963 2117 1966
rect 2082 1913 2085 1936
rect 2082 1803 2085 1906
rect 2090 1853 2093 1925
rect 2098 1923 2101 1963
rect 2122 1956 2125 1976
rect 2106 1933 2109 1956
rect 2114 1953 2125 1956
rect 2106 1906 2109 1926
rect 2098 1903 2109 1906
rect 2098 1873 2101 1903
rect 2090 1823 2101 1826
rect 2090 1796 2093 1823
rect 2082 1793 2093 1796
rect 2058 1503 2061 1516
rect 2058 1376 2061 1466
rect 2066 1393 2069 1523
rect 2074 1483 2077 1516
rect 2074 1383 2077 1416
rect 2082 1393 2085 1793
rect 2098 1766 2101 1816
rect 2106 1813 2109 1896
rect 2114 1803 2117 1953
rect 2122 1913 2125 1926
rect 2122 1773 2125 1896
rect 2098 1763 2125 1766
rect 2090 1526 2093 1726
rect 2098 1636 2101 1763
rect 2106 1733 2109 1746
rect 2106 1696 2109 1726
rect 2114 1716 2117 1756
rect 2122 1733 2125 1763
rect 2114 1713 2125 1716
rect 2130 1696 2133 2166
rect 2146 2143 2149 2186
rect 2138 2013 2141 2036
rect 2138 1923 2141 1936
rect 2138 1823 2141 1916
rect 2146 1893 2149 2086
rect 2146 1816 2149 1826
rect 2154 1823 2157 2256
rect 2162 2036 2165 2343
rect 2178 2333 2181 2416
rect 2218 2413 2221 2426
rect 2202 2333 2205 2356
rect 2186 2323 2197 2326
rect 2202 2323 2213 2326
rect 2178 2266 2181 2316
rect 2178 2263 2189 2266
rect 2170 2156 2173 2216
rect 2178 2213 2181 2256
rect 2170 2153 2181 2156
rect 2170 2133 2173 2146
rect 2170 2103 2173 2126
rect 2178 2073 2181 2153
rect 2162 2033 2173 2036
rect 2162 2013 2165 2026
rect 2162 1953 2165 2006
rect 2170 1936 2173 2033
rect 2178 2023 2181 2046
rect 2162 1933 2173 1936
rect 2162 1913 2165 1933
rect 2170 1873 2173 1926
rect 2138 1813 2149 1816
rect 2138 1736 2141 1813
rect 2146 1753 2149 1806
rect 2138 1733 2149 1736
rect 2154 1733 2157 1816
rect 2162 1766 2165 1806
rect 2178 1773 2181 1936
rect 2186 1916 2189 2263
rect 2194 2206 2197 2226
rect 2202 2213 2205 2323
rect 2226 2273 2229 2443
rect 2234 2423 2237 2526
rect 2266 2523 2269 2556
rect 2242 2376 2245 2416
rect 2266 2383 2269 2426
rect 2274 2413 2277 2573
rect 2282 2483 2285 2616
rect 2298 2533 2301 2616
rect 2314 2613 2317 2696
rect 2322 2546 2325 2626
rect 2338 2603 2341 2616
rect 2362 2576 2365 2646
rect 2378 2606 2381 2776
rect 2450 2766 2453 2816
rect 2458 2796 2461 2823
rect 2458 2793 2469 2796
rect 2458 2773 2461 2786
rect 2418 2763 2453 2766
rect 2386 2733 2389 2756
rect 2410 2716 2413 2726
rect 2418 2723 2421 2763
rect 2410 2713 2421 2716
rect 2410 2686 2413 2706
rect 2406 2683 2413 2686
rect 2338 2573 2365 2576
rect 2370 2603 2381 2606
rect 2322 2543 2329 2546
rect 2274 2376 2277 2406
rect 2242 2373 2277 2376
rect 2282 2353 2285 2446
rect 2298 2403 2301 2526
rect 2326 2496 2329 2543
rect 2322 2493 2329 2496
rect 2306 2393 2309 2406
rect 2314 2403 2317 2426
rect 2322 2343 2325 2493
rect 2338 2436 2341 2573
rect 2346 2486 2349 2526
rect 2370 2493 2373 2603
rect 2378 2523 2381 2596
rect 2386 2566 2389 2616
rect 2386 2563 2393 2566
rect 2346 2483 2381 2486
rect 2334 2433 2341 2436
rect 2334 2356 2337 2433
rect 2334 2353 2341 2356
rect 2338 2336 2341 2353
rect 2242 2306 2245 2336
rect 2258 2333 2341 2336
rect 2258 2313 2261 2333
rect 2242 2303 2261 2306
rect 2210 2216 2213 2236
rect 2218 2223 2221 2266
rect 2234 2226 2237 2236
rect 2226 2223 2237 2226
rect 2226 2216 2229 2223
rect 2210 2213 2229 2216
rect 2234 2206 2237 2216
rect 2242 2213 2245 2303
rect 2194 2203 2237 2206
rect 2234 2193 2237 2203
rect 2194 2103 2197 2126
rect 2202 2023 2205 2136
rect 2218 2123 2221 2166
rect 2234 2133 2245 2136
rect 2210 2093 2213 2106
rect 2218 2083 2221 2116
rect 2234 2113 2237 2133
rect 2250 2076 2253 2296
rect 2258 2223 2261 2236
rect 2266 2223 2269 2326
rect 2274 2313 2301 2316
rect 2258 2083 2261 2146
rect 2266 2076 2269 2176
rect 2226 2073 2253 2076
rect 2258 2073 2269 2076
rect 2226 2056 2229 2073
rect 2222 2053 2229 2056
rect 2194 1973 2197 2006
rect 2202 1993 2205 2006
rect 2222 1996 2225 2053
rect 2210 1956 2213 1996
rect 2218 1993 2225 1996
rect 2218 1976 2221 1993
rect 2234 1986 2237 2036
rect 2226 1983 2237 1986
rect 2242 1983 2245 2006
rect 2250 2003 2253 2016
rect 2258 1996 2261 2073
rect 2250 1993 2261 1996
rect 2266 1993 2269 2066
rect 2274 2013 2277 2313
rect 2282 2063 2285 2266
rect 2290 2233 2293 2306
rect 2306 2236 2309 2326
rect 2298 2233 2309 2236
rect 2290 2026 2293 2146
rect 2282 2023 2293 2026
rect 2298 2023 2301 2226
rect 2306 2213 2309 2226
rect 2314 2196 2317 2276
rect 2322 2233 2325 2326
rect 2310 2193 2317 2196
rect 2310 2116 2313 2193
rect 2322 2133 2325 2186
rect 2330 2163 2333 2316
rect 2338 2233 2341 2333
rect 2346 2273 2349 2426
rect 2354 2403 2357 2426
rect 2362 2416 2365 2476
rect 2378 2416 2381 2483
rect 2390 2446 2393 2563
rect 2406 2556 2409 2683
rect 2418 2613 2421 2713
rect 2442 2686 2445 2736
rect 2466 2723 2469 2793
rect 2474 2766 2477 2856
rect 2490 2853 2533 2856
rect 2490 2813 2493 2853
rect 2530 2813 2533 2853
rect 2546 2836 2549 2883
rect 2566 2866 2569 2963
rect 2590 2906 2593 2993
rect 2586 2903 2593 2906
rect 2586 2886 2589 2903
rect 2578 2883 2589 2886
rect 2566 2863 2573 2866
rect 2546 2833 2557 2836
rect 2554 2813 2557 2833
rect 2506 2793 2509 2806
rect 2570 2773 2573 2863
rect 2578 2766 2581 2883
rect 2602 2816 2605 2926
rect 2610 2923 2613 2946
rect 2618 2933 2621 3016
rect 2626 3013 2629 3023
rect 2634 3016 2637 3143
rect 2642 3133 2653 3136
rect 2658 3126 2661 3213
rect 2666 3143 2669 3216
rect 2714 3203 2717 3226
rect 2794 3216 2797 3236
rect 2738 3193 2741 3216
rect 2786 3213 2797 3216
rect 2682 3133 2685 3146
rect 2690 3143 2733 3146
rect 2690 3133 2693 3143
rect 2714 3133 2725 3136
rect 2730 3133 2733 3143
rect 2738 3133 2741 3166
rect 2642 3123 2661 3126
rect 2666 3123 2757 3126
rect 2642 3103 2645 3123
rect 2658 3083 2661 3116
rect 2634 3013 2653 3016
rect 2626 2993 2629 3006
rect 2642 3003 2653 3006
rect 2642 2946 2645 3003
rect 2666 2996 2669 3016
rect 2674 3013 2677 3026
rect 2682 3013 2685 3026
rect 2690 3006 2693 3056
rect 2650 2993 2669 2996
rect 2674 3003 2693 3006
rect 2642 2943 2669 2946
rect 2626 2933 2637 2936
rect 2666 2933 2669 2943
rect 2626 2923 2637 2926
rect 2626 2893 2629 2923
rect 2666 2916 2669 2926
rect 2634 2913 2669 2916
rect 2474 2763 2525 2766
rect 2522 2723 2525 2763
rect 2562 2763 2581 2766
rect 2530 2733 2533 2746
rect 2546 2713 2549 2726
rect 2562 2723 2565 2763
rect 2570 2733 2573 2756
rect 2578 2696 2581 2763
rect 2586 2723 2589 2816
rect 2602 2813 2621 2816
rect 2626 2806 2629 2846
rect 2634 2813 2637 2826
rect 2674 2816 2677 3003
rect 2706 2986 2709 3116
rect 2762 3083 2765 3136
rect 2786 3123 2789 3213
rect 2802 3106 2805 3126
rect 2794 3103 2805 3106
rect 2714 3033 2749 3036
rect 2714 2993 2717 3033
rect 2746 3013 2749 3033
rect 2722 2986 2725 3006
rect 2706 2983 2725 2986
rect 2682 2923 2685 2936
rect 2690 2933 2693 2956
rect 2770 2943 2773 3006
rect 2722 2933 2773 2936
rect 2778 2926 2781 3016
rect 2794 2966 2797 3103
rect 2810 3036 2813 3136
rect 2802 3033 2813 3036
rect 2802 3003 2805 3033
rect 2818 2976 2821 3176
rect 2826 3123 2829 3206
rect 2842 3113 2845 3146
rect 2850 3133 2853 3216
rect 2818 2973 2837 2976
rect 2794 2963 2829 2966
rect 2722 2913 2725 2926
rect 2730 2843 2733 2926
rect 2746 2836 2749 2926
rect 2754 2923 2781 2926
rect 2754 2913 2757 2923
rect 2746 2833 2753 2836
rect 2602 2773 2605 2806
rect 2610 2803 2629 2806
rect 2578 2693 2589 2696
rect 2442 2683 2477 2686
rect 2418 2586 2421 2606
rect 2442 2603 2445 2616
rect 2418 2583 2425 2586
rect 2406 2553 2413 2556
rect 2386 2443 2393 2446
rect 2386 2423 2389 2443
rect 2362 2413 2373 2416
rect 2378 2413 2389 2416
rect 2362 2393 2365 2406
rect 2370 2363 2373 2413
rect 2386 2403 2389 2413
rect 2338 2193 2341 2226
rect 2346 2206 2349 2246
rect 2354 2223 2357 2326
rect 2362 2213 2365 2226
rect 2346 2203 2353 2206
rect 2338 2126 2341 2146
rect 2350 2136 2353 2203
rect 2370 2176 2373 2346
rect 2378 2323 2389 2326
rect 2394 2313 2397 2426
rect 2402 2393 2405 2536
rect 2402 2333 2405 2376
rect 2410 2333 2413 2553
rect 2422 2506 2425 2583
rect 2466 2576 2469 2616
rect 2434 2573 2469 2576
rect 2434 2533 2437 2573
rect 2474 2566 2477 2683
rect 2522 2613 2525 2656
rect 2586 2626 2589 2693
rect 2610 2673 2613 2803
rect 2582 2623 2589 2626
rect 2450 2563 2477 2566
rect 2450 2533 2453 2563
rect 2474 2546 2477 2563
rect 2474 2543 2485 2546
rect 2418 2503 2425 2506
rect 2402 2323 2413 2326
rect 2362 2173 2373 2176
rect 2362 2153 2365 2173
rect 2350 2133 2357 2136
rect 2322 2123 2341 2126
rect 2310 2113 2317 2116
rect 2218 1973 2245 1976
rect 2194 1953 2213 1956
rect 2194 1943 2197 1953
rect 2226 1946 2229 1956
rect 2210 1943 2229 1946
rect 2210 1923 2213 1936
rect 2186 1913 2197 1916
rect 2162 1763 2181 1766
rect 2138 1703 2141 1726
rect 2106 1693 2117 1696
rect 2130 1693 2141 1696
rect 2106 1656 2109 1686
rect 2114 1663 2117 1693
rect 2106 1653 2133 1656
rect 2098 1633 2125 1636
rect 2130 1626 2133 1653
rect 2122 1623 2133 1626
rect 2098 1603 2101 1616
rect 2098 1556 2101 1586
rect 2106 1563 2109 1606
rect 2114 1603 2117 1616
rect 2122 1596 2125 1623
rect 2122 1593 2133 1596
rect 2098 1553 2109 1556
rect 2090 1523 2101 1526
rect 2098 1503 2101 1523
rect 2058 1373 2065 1376
rect 2062 1246 2065 1373
rect 2074 1293 2077 1326
rect 2082 1303 2085 1336
rect 2058 1243 2065 1246
rect 2058 1093 2061 1243
rect 2066 1133 2069 1226
rect 2082 1133 2085 1216
rect 2090 1153 2093 1466
rect 2098 1283 2101 1496
rect 2106 1463 2109 1553
rect 2114 1533 2117 1556
rect 2122 1533 2125 1566
rect 2130 1526 2133 1593
rect 2122 1523 2133 1526
rect 2058 963 2061 1016
rect 2066 1006 2069 1106
rect 2074 1013 2077 1126
rect 2090 1113 2093 1126
rect 2098 1123 2101 1186
rect 2082 1103 2101 1106
rect 2082 1073 2085 1103
rect 2098 1076 2101 1096
rect 2094 1073 2101 1076
rect 2066 1003 2077 1006
rect 2050 943 2057 946
rect 2054 836 2057 943
rect 2066 933 2069 996
rect 2074 923 2077 986
rect 2082 923 2085 1016
rect 2094 1006 2097 1073
rect 2106 1023 2109 1426
rect 2094 1003 2101 1006
rect 2098 986 2101 1003
rect 2106 993 2109 1016
rect 2098 983 2109 986
rect 2050 833 2057 836
rect 2002 823 2029 826
rect 1994 706 1997 816
rect 2002 786 2005 823
rect 2010 803 2013 816
rect 2002 783 2009 786
rect 1986 703 1997 706
rect 1986 646 1989 703
rect 2006 696 2009 783
rect 2002 693 2009 696
rect 1986 643 1997 646
rect 1970 623 1981 626
rect 1946 593 1957 596
rect 1962 596 1965 616
rect 1962 593 1969 596
rect 1946 576 1949 593
rect 1942 573 1949 576
rect 1898 503 1901 516
rect 1878 423 1885 426
rect 1858 393 1869 396
rect 1866 316 1869 393
rect 1878 326 1881 423
rect 1890 333 1893 416
rect 1898 333 1901 496
rect 1878 323 1885 326
rect 1906 323 1909 533
rect 1914 523 1925 526
rect 1930 436 1933 536
rect 1942 516 1945 573
rect 1954 523 1957 566
rect 1942 513 1949 516
rect 1914 433 1933 436
rect 1914 423 1917 433
rect 1922 423 1933 426
rect 1914 373 1917 406
rect 1922 376 1925 416
rect 1946 413 1949 513
rect 1966 496 1969 593
rect 1962 493 1969 496
rect 1962 473 1965 493
rect 1978 466 1981 623
rect 1994 593 1997 643
rect 2002 586 2005 693
rect 2010 613 2013 636
rect 1994 583 2005 586
rect 1994 526 1997 583
rect 2010 563 2013 606
rect 2018 593 2021 816
rect 2042 813 2045 826
rect 2026 803 2037 806
rect 2042 793 2045 806
rect 2050 776 2053 833
rect 2034 733 2037 776
rect 2046 773 2053 776
rect 2026 706 2029 726
rect 2046 716 2049 773
rect 2058 723 2061 816
rect 2066 793 2069 856
rect 2074 786 2077 906
rect 2070 783 2077 786
rect 2070 716 2073 783
rect 2046 713 2053 716
rect 2026 703 2037 706
rect 2034 646 2037 703
rect 2026 643 2037 646
rect 2026 626 2029 643
rect 2026 623 2037 626
rect 1970 463 1981 466
rect 1990 523 1997 526
rect 1990 466 1993 523
rect 2002 476 2005 536
rect 2026 533 2029 576
rect 2042 533 2045 626
rect 2050 586 2053 713
rect 2066 713 2073 716
rect 2058 603 2061 646
rect 2050 583 2057 586
rect 2010 523 2029 526
rect 2026 486 2029 516
rect 2026 483 2037 486
rect 2002 473 2029 476
rect 1990 463 1997 466
rect 1930 383 1933 406
rect 1970 383 1973 463
rect 1922 373 1941 376
rect 1834 313 1853 316
rect 1858 313 1869 316
rect 1802 273 1813 276
rect 1778 163 1797 166
rect 1746 116 1749 146
rect 1754 143 1765 146
rect 1738 113 1749 116
rect 1634 83 1645 86
rect 1738 36 1741 113
rect 1762 56 1765 143
rect 1786 123 1789 146
rect 1794 116 1797 163
rect 1802 123 1805 266
rect 1810 123 1813 273
rect 1818 123 1821 216
rect 1834 203 1837 313
rect 1858 293 1861 313
rect 1850 223 1853 236
rect 1850 176 1853 206
rect 1826 173 1853 176
rect 1826 123 1829 166
rect 1882 163 1885 323
rect 1922 306 1925 336
rect 1930 313 1933 346
rect 1938 333 1941 373
rect 1978 366 1981 416
rect 1994 386 1997 463
rect 2026 413 2029 473
rect 2034 463 2037 483
rect 2010 403 2021 406
rect 2034 403 2037 436
rect 2042 423 2045 516
rect 2054 436 2057 583
rect 2050 433 2057 436
rect 2002 393 2013 396
rect 1970 363 1981 366
rect 1970 316 1973 363
rect 1914 303 1925 306
rect 1914 216 1917 303
rect 1914 213 1925 216
rect 1922 196 1925 213
rect 1890 193 1925 196
rect 1930 193 1933 206
rect 1938 166 1941 316
rect 1970 313 1981 316
rect 1978 223 1981 313
rect 1946 173 1949 216
rect 1986 203 1989 386
rect 1994 383 2013 386
rect 1994 286 1997 316
rect 2002 306 2005 326
rect 2010 323 2013 383
rect 2018 333 2021 403
rect 2042 373 2045 416
rect 2026 323 2029 366
rect 2034 306 2037 336
rect 2002 303 2037 306
rect 1994 283 2005 286
rect 2002 236 2005 283
rect 2050 276 2053 433
rect 2066 426 2069 713
rect 2074 493 2077 626
rect 2066 423 2073 426
rect 2058 383 2061 416
rect 2070 366 2073 423
rect 2082 373 2085 856
rect 2090 633 2093 976
rect 2098 903 2101 966
rect 2106 853 2109 983
rect 2114 963 2117 1516
rect 2122 1366 2125 1523
rect 2138 1503 2141 1693
rect 2146 1563 2149 1733
rect 2154 1713 2157 1726
rect 2154 1623 2157 1636
rect 2138 1483 2141 1496
rect 2130 1383 2133 1456
rect 2138 1403 2141 1476
rect 2146 1423 2149 1536
rect 2154 1533 2157 1606
rect 2154 1416 2157 1516
rect 2162 1496 2165 1756
rect 2170 1733 2173 1746
rect 2178 1726 2181 1763
rect 2186 1743 2189 1886
rect 2194 1803 2197 1913
rect 2218 1906 2221 1936
rect 2214 1903 2221 1906
rect 2194 1733 2197 1796
rect 2170 1653 2173 1726
rect 2178 1723 2185 1726
rect 2182 1616 2185 1723
rect 2194 1653 2197 1726
rect 2202 1676 2205 1846
rect 2214 1836 2217 1903
rect 2226 1863 2229 1943
rect 2210 1833 2217 1836
rect 2210 1793 2213 1833
rect 2234 1826 2237 1936
rect 2242 1933 2245 1973
rect 2250 1933 2253 1993
rect 2242 1843 2245 1926
rect 2258 1893 2261 1986
rect 2266 1923 2269 1976
rect 2274 1933 2277 2006
rect 2282 1986 2285 2023
rect 2290 2003 2293 2016
rect 2298 1993 2301 2006
rect 2282 1983 2289 1986
rect 2218 1823 2237 1826
rect 2210 1683 2213 1786
rect 2202 1673 2213 1676
rect 2194 1623 2197 1646
rect 2182 1613 2189 1616
rect 2170 1523 2173 1556
rect 2178 1513 2181 1606
rect 2186 1603 2189 1613
rect 2186 1523 2189 1546
rect 2194 1506 2197 1606
rect 2202 1523 2205 1616
rect 2210 1603 2213 1673
rect 2210 1543 2213 1566
rect 2190 1503 2197 1506
rect 2162 1493 2173 1496
rect 2170 1426 2173 1493
rect 2190 1446 2193 1503
rect 2190 1443 2197 1446
rect 2170 1423 2189 1426
rect 2122 1363 2129 1366
rect 2126 1156 2129 1363
rect 2122 1153 2129 1156
rect 2122 1093 2125 1153
rect 2130 1016 2133 1136
rect 2122 1013 2133 1016
rect 2122 933 2125 1013
rect 2130 916 2133 1006
rect 2138 993 2141 1396
rect 2146 1333 2149 1416
rect 2154 1413 2165 1416
rect 2154 1373 2157 1406
rect 2162 1336 2165 1413
rect 2178 1393 2181 1416
rect 2154 1333 2165 1336
rect 2170 1333 2173 1346
rect 2146 943 2149 1216
rect 2154 1173 2157 1333
rect 2162 1323 2173 1326
rect 2170 1223 2173 1323
rect 2170 1153 2173 1186
rect 2178 1136 2181 1386
rect 2154 1113 2157 1136
rect 2170 1133 2181 1136
rect 2186 1133 2189 1423
rect 2170 1113 2173 1133
rect 2194 1126 2197 1443
rect 2202 1403 2205 1516
rect 2202 1233 2205 1326
rect 2210 1233 2213 1536
rect 2202 1203 2205 1226
rect 2210 1173 2213 1206
rect 2178 1123 2197 1126
rect 2154 1003 2157 1076
rect 2114 913 2133 916
rect 2098 803 2101 826
rect 2114 823 2117 913
rect 2098 743 2117 746
rect 2098 733 2109 736
rect 2090 433 2093 626
rect 2098 513 2101 706
rect 2106 603 2109 733
rect 2114 686 2117 736
rect 2122 703 2125 906
rect 2130 803 2133 906
rect 2138 806 2141 926
rect 2146 923 2157 926
rect 2154 903 2157 916
rect 2162 863 2165 936
rect 2146 813 2149 856
rect 2138 803 2149 806
rect 2130 793 2141 796
rect 2130 743 2133 793
rect 2114 683 2121 686
rect 2118 596 2121 683
rect 2114 593 2121 596
rect 2114 526 2117 593
rect 2130 533 2133 646
rect 2138 593 2141 756
rect 2106 523 2117 526
rect 2130 523 2141 526
rect 2066 363 2073 366
rect 2066 333 2069 363
rect 2074 316 2077 346
rect 2098 336 2101 496
rect 2106 433 2109 523
rect 2130 516 2133 523
rect 2114 513 2133 516
rect 2146 506 2149 803
rect 2154 803 2165 806
rect 2154 733 2157 803
rect 2170 793 2173 966
rect 2178 906 2181 1123
rect 2186 923 2189 1006
rect 2178 903 2185 906
rect 2182 836 2185 903
rect 2178 833 2185 836
rect 2178 813 2181 833
rect 2194 816 2197 1076
rect 2202 1026 2205 1166
rect 2218 1073 2221 1823
rect 2242 1816 2245 1826
rect 2250 1823 2253 1886
rect 2274 1856 2277 1926
rect 2286 1896 2289 1983
rect 2306 1956 2309 2016
rect 2314 1973 2317 2113
rect 2338 2106 2341 2123
rect 2334 2103 2341 2106
rect 2334 2036 2337 2103
rect 2346 2043 2349 2126
rect 2354 2093 2357 2133
rect 2370 2123 2373 2166
rect 2378 2156 2381 2226
rect 2386 2223 2389 2266
rect 2394 2233 2397 2286
rect 2418 2276 2421 2503
rect 2426 2416 2429 2486
rect 2434 2443 2437 2516
rect 2482 2496 2485 2543
rect 2498 2523 2501 2536
rect 2554 2533 2557 2616
rect 2434 2423 2445 2426
rect 2426 2413 2437 2416
rect 2434 2403 2437 2413
rect 2426 2316 2429 2386
rect 2434 2333 2437 2396
rect 2442 2373 2445 2406
rect 2450 2393 2453 2496
rect 2474 2493 2485 2496
rect 2474 2436 2477 2493
rect 2474 2433 2501 2436
rect 2466 2403 2469 2416
rect 2474 2396 2477 2433
rect 2466 2393 2477 2396
rect 2466 2333 2469 2393
rect 2482 2373 2485 2426
rect 2498 2403 2501 2433
rect 2538 2426 2541 2526
rect 2582 2436 2585 2623
rect 2594 2476 2597 2616
rect 2634 2613 2637 2716
rect 2642 2596 2645 2816
rect 2658 2813 2685 2816
rect 2650 2743 2653 2806
rect 2674 2753 2677 2806
rect 2682 2736 2685 2813
rect 2698 2803 2701 2816
rect 2738 2813 2741 2826
rect 2714 2793 2717 2806
rect 2750 2766 2753 2833
rect 2794 2803 2797 2816
rect 2802 2796 2805 2946
rect 2826 2923 2829 2963
rect 2834 2843 2837 2973
rect 2858 2966 2861 3166
rect 2866 3013 2869 3026
rect 2850 2963 2861 2966
rect 2818 2803 2821 2826
rect 2826 2813 2829 2836
rect 2786 2793 2805 2796
rect 2750 2763 2757 2766
rect 2678 2733 2685 2736
rect 2658 2693 2661 2726
rect 2650 2603 2653 2676
rect 2678 2636 2681 2733
rect 2690 2643 2693 2726
rect 2678 2633 2685 2636
rect 2682 2613 2685 2633
rect 2634 2593 2645 2596
rect 2634 2546 2637 2593
rect 2602 2523 2605 2546
rect 2634 2543 2645 2546
rect 2642 2523 2645 2543
rect 2642 2496 2645 2516
rect 2650 2503 2653 2536
rect 2634 2493 2645 2496
rect 2594 2473 2605 2476
rect 2582 2433 2589 2436
rect 2530 2423 2541 2426
rect 2530 2376 2533 2423
rect 2586 2416 2589 2433
rect 2602 2416 2605 2473
rect 2634 2446 2637 2493
rect 2658 2446 2661 2586
rect 2698 2556 2701 2606
rect 2706 2603 2709 2616
rect 2714 2596 2717 2736
rect 2722 2703 2725 2726
rect 2738 2673 2741 2716
rect 2754 2666 2757 2763
rect 2730 2663 2757 2666
rect 2730 2646 2733 2663
rect 2706 2593 2717 2596
rect 2726 2643 2733 2646
rect 2726 2566 2729 2643
rect 2738 2613 2741 2636
rect 2746 2613 2749 2626
rect 2726 2563 2733 2566
rect 2682 2553 2701 2556
rect 2674 2533 2677 2546
rect 2634 2443 2645 2446
rect 2658 2443 2669 2446
rect 2530 2373 2541 2376
rect 2490 2346 2493 2366
rect 2490 2343 2501 2346
rect 2426 2313 2437 2316
rect 2410 2273 2421 2276
rect 2410 2233 2413 2273
rect 2418 2233 2421 2266
rect 2434 2236 2437 2313
rect 2426 2233 2437 2236
rect 2394 2213 2397 2226
rect 2410 2163 2413 2226
rect 2418 2213 2421 2226
rect 2378 2153 2389 2156
rect 2378 2133 2381 2146
rect 2378 2113 2381 2126
rect 2334 2033 2341 2036
rect 2322 1993 2325 2026
rect 2338 2016 2341 2033
rect 2362 2016 2365 2026
rect 2298 1953 2309 1956
rect 2298 1943 2301 1953
rect 2314 1946 2317 1966
rect 2306 1943 2317 1946
rect 2298 1923 2301 1936
rect 2314 1926 2317 1943
rect 2310 1923 2317 1926
rect 2322 1923 2325 1936
rect 2286 1893 2293 1896
rect 2266 1853 2277 1856
rect 2226 1773 2229 1806
rect 2234 1796 2237 1816
rect 2242 1813 2253 1816
rect 2258 1813 2261 1826
rect 2250 1803 2253 1813
rect 2234 1793 2253 1796
rect 2226 1733 2245 1736
rect 2250 1733 2253 1793
rect 2258 1783 2261 1806
rect 2226 1723 2229 1733
rect 2242 1726 2245 1733
rect 2234 1706 2237 1726
rect 2242 1723 2253 1726
rect 2226 1703 2237 1706
rect 2250 1686 2253 1716
rect 2258 1713 2261 1766
rect 2266 1686 2269 1853
rect 2274 1813 2277 1846
rect 2282 1823 2285 1886
rect 2290 1843 2293 1893
rect 2274 1803 2285 1806
rect 2290 1733 2293 1826
rect 2298 1823 2301 1916
rect 2310 1846 2313 1923
rect 2330 1876 2333 2016
rect 2338 2013 2365 2016
rect 2338 1963 2341 2013
rect 2354 1946 2357 2006
rect 2370 1993 2373 2066
rect 2386 2053 2389 2153
rect 2394 2133 2405 2136
rect 2410 2133 2413 2146
rect 2402 2113 2405 2126
rect 2378 1956 2381 2046
rect 2386 2013 2389 2026
rect 2338 1933 2341 1946
rect 2346 1943 2357 1946
rect 2362 1953 2381 1956
rect 2330 1873 2337 1876
rect 2306 1843 2313 1846
rect 2298 1793 2301 1816
rect 2306 1803 2309 1843
rect 2274 1703 2277 1726
rect 2282 1723 2293 1726
rect 2298 1716 2301 1746
rect 2314 1716 2317 1826
rect 2322 1763 2325 1866
rect 2334 1816 2337 1873
rect 2346 1863 2349 1943
rect 2354 1853 2357 1936
rect 2362 1923 2365 1953
rect 2386 1936 2389 1996
rect 2394 1966 2397 2006
rect 2402 1993 2405 2056
rect 2410 1993 2413 2076
rect 2418 1993 2421 2156
rect 2394 1963 2405 1966
rect 2394 1943 2397 1956
rect 2370 1913 2373 1936
rect 2386 1933 2397 1936
rect 2346 1816 2349 1836
rect 2354 1823 2365 1826
rect 2334 1813 2341 1816
rect 2346 1813 2357 1816
rect 2330 1793 2333 1806
rect 2290 1713 2301 1716
rect 2310 1713 2317 1716
rect 2250 1683 2261 1686
rect 2266 1683 2285 1686
rect 2226 1623 2229 1666
rect 2258 1656 2261 1683
rect 2226 1553 2229 1616
rect 2242 1556 2245 1636
rect 2234 1553 2245 1556
rect 2226 1506 2229 1526
rect 2234 1523 2237 1553
rect 2250 1533 2253 1656
rect 2258 1653 2269 1656
rect 2266 1613 2269 1653
rect 2282 1643 2285 1683
rect 2274 1613 2285 1616
rect 2258 1583 2261 1606
rect 2282 1543 2285 1606
rect 2290 1526 2293 1713
rect 2298 1606 2301 1686
rect 2310 1656 2313 1713
rect 2310 1653 2317 1656
rect 2306 1613 2309 1636
rect 2298 1603 2309 1606
rect 2298 1533 2301 1596
rect 2226 1503 2233 1506
rect 2230 1436 2233 1503
rect 2226 1433 2233 1436
rect 2226 1413 2229 1433
rect 2242 1423 2245 1526
rect 2226 1333 2229 1406
rect 2258 1353 2261 1416
rect 2242 1323 2245 1336
rect 2226 1133 2229 1266
rect 2234 1213 2237 1276
rect 2242 1213 2245 1226
rect 2250 1193 2253 1346
rect 2266 1196 2269 1526
rect 2282 1523 2293 1526
rect 2282 1456 2285 1523
rect 2282 1453 2293 1456
rect 2282 1413 2285 1436
rect 2274 1403 2285 1406
rect 2290 1383 2293 1453
rect 2298 1413 2301 1526
rect 2306 1513 2309 1603
rect 2282 1333 2301 1336
rect 2274 1306 2277 1326
rect 2298 1323 2301 1333
rect 2274 1303 2285 1306
rect 2298 1303 2301 1316
rect 2282 1236 2285 1303
rect 2274 1233 2285 1236
rect 2274 1203 2277 1233
rect 2298 1223 2301 1256
rect 2282 1213 2301 1216
rect 2266 1193 2285 1196
rect 2210 1033 2221 1036
rect 2202 1023 2209 1026
rect 2206 966 2209 1023
rect 2206 963 2213 966
rect 2202 933 2205 946
rect 2210 816 2213 963
rect 2218 943 2221 1033
rect 2226 1013 2229 1126
rect 2234 1106 2237 1166
rect 2242 1123 2245 1186
rect 2250 1133 2277 1136
rect 2250 1116 2253 1133
rect 2242 1113 2253 1116
rect 2258 1123 2269 1126
rect 2274 1123 2277 1133
rect 2234 1103 2241 1106
rect 2238 1036 2241 1103
rect 2238 1033 2245 1036
rect 2234 1003 2237 1016
rect 2218 903 2221 936
rect 2226 843 2229 926
rect 2242 826 2245 1033
rect 2250 923 2253 1096
rect 2258 1013 2261 1123
rect 2282 1116 2285 1193
rect 2274 1113 2285 1116
rect 2242 823 2253 826
rect 2190 813 2197 816
rect 2202 813 2221 816
rect 2190 756 2193 813
rect 2162 723 2165 756
rect 2190 753 2197 756
rect 2186 716 2189 736
rect 2194 733 2197 753
rect 2154 516 2157 686
rect 2162 533 2165 616
rect 2170 566 2173 656
rect 2178 596 2181 716
rect 2186 713 2193 716
rect 2190 636 2193 713
rect 2186 633 2193 636
rect 2186 606 2189 633
rect 2202 623 2205 813
rect 2218 796 2221 806
rect 2210 793 2221 796
rect 2210 753 2213 793
rect 2218 766 2221 786
rect 2234 776 2237 806
rect 2226 773 2237 776
rect 2242 773 2245 796
rect 2218 763 2229 766
rect 2226 673 2229 763
rect 2210 623 2229 626
rect 2194 613 2205 616
rect 2186 603 2197 606
rect 2178 593 2189 596
rect 2170 563 2181 566
rect 2154 513 2161 516
rect 2138 503 2149 506
rect 2114 373 2117 416
rect 2130 373 2133 426
rect 2138 346 2141 503
rect 2146 406 2149 496
rect 2158 446 2161 513
rect 2170 493 2173 546
rect 2178 533 2181 563
rect 2186 483 2189 593
rect 2154 443 2161 446
rect 2154 416 2157 443
rect 2162 423 2189 426
rect 2194 423 2197 603
rect 2202 543 2205 613
rect 2202 433 2205 526
rect 2154 413 2181 416
rect 2146 403 2157 406
rect 2134 343 2141 346
rect 2082 333 2101 336
rect 2082 323 2085 333
rect 2074 313 2085 316
rect 2082 296 2085 313
rect 2098 306 2101 326
rect 2106 313 2109 336
rect 2098 303 2109 306
rect 2082 293 2089 296
rect 1994 233 2005 236
rect 2042 273 2053 276
rect 1994 213 1997 233
rect 2042 226 2045 273
rect 2042 223 2053 226
rect 2034 196 2037 206
rect 1954 193 2037 196
rect 1938 163 1965 166
rect 1834 116 1837 126
rect 1794 113 1837 116
rect 1898 103 1901 136
rect 1922 133 1925 146
rect 1906 83 1909 126
rect 1954 116 1957 136
rect 1962 123 1965 163
rect 1970 116 1973 136
rect 1754 53 1765 56
rect 1738 33 1749 36
rect 1754 33 1757 53
rect 1922 43 1925 116
rect 1954 113 1973 116
rect 1978 53 1981 126
rect 1986 43 1989 166
rect 1746 13 1749 33
rect 2034 23 2037 136
rect 2042 123 2045 206
rect 2050 133 2053 223
rect 2058 133 2061 266
rect 2066 143 2069 226
rect 2074 213 2077 266
rect 2086 206 2089 293
rect 2098 213 2101 303
rect 2114 293 2117 326
rect 2134 286 2137 343
rect 2146 293 2149 316
rect 2154 313 2157 403
rect 2170 326 2173 406
rect 2178 363 2181 413
rect 2186 333 2189 423
rect 2170 323 2189 326
rect 2194 313 2197 416
rect 2202 393 2205 406
rect 2210 313 2213 623
rect 2170 296 2173 306
rect 2218 296 2221 616
rect 2226 613 2229 623
rect 2242 606 2245 726
rect 2250 686 2253 823
rect 2258 703 2261 986
rect 2266 933 2269 1026
rect 2274 916 2277 1113
rect 2282 1023 2285 1076
rect 2270 913 2277 916
rect 2270 806 2273 913
rect 2282 823 2285 936
rect 2270 803 2277 806
rect 2274 783 2277 803
rect 2266 743 2269 776
rect 2282 726 2285 816
rect 2290 783 2293 1126
rect 2274 723 2285 726
rect 2250 683 2261 686
rect 2258 636 2261 683
rect 2250 633 2261 636
rect 2250 613 2253 633
rect 2274 626 2277 723
rect 2290 706 2293 736
rect 2286 703 2293 706
rect 2286 646 2289 703
rect 2298 653 2301 1206
rect 2306 1133 2309 1416
rect 2306 943 2309 1126
rect 2306 863 2309 916
rect 2306 683 2309 836
rect 2286 643 2293 646
rect 2274 623 2285 626
rect 2226 583 2229 606
rect 2242 603 2277 606
rect 2226 533 2229 546
rect 2170 293 2189 296
rect 2134 283 2141 286
rect 2106 213 2109 276
rect 2082 203 2089 206
rect 2122 203 2125 226
rect 2058 113 2061 126
rect 2082 123 2085 203
rect 2114 46 2117 136
rect 2130 133 2133 166
rect 2138 113 2141 283
rect 2162 213 2165 276
rect 2186 236 2189 293
rect 2178 233 2189 236
rect 2210 293 2221 296
rect 2178 213 2181 233
rect 2210 226 2213 293
rect 2210 223 2221 226
rect 2146 53 2149 136
rect 2162 126 2165 136
rect 2154 46 2157 126
rect 2162 123 2181 126
rect 2162 106 2165 123
rect 2162 103 2173 106
rect 2170 46 2173 103
rect 2114 43 2157 46
rect 2162 43 2173 46
rect 2162 23 2165 43
rect 2186 33 2189 216
rect 2194 176 2197 206
rect 2218 193 2221 223
rect 2226 213 2229 516
rect 2234 423 2237 596
rect 2234 313 2237 376
rect 2242 213 2245 603
rect 2250 593 2261 596
rect 2274 593 2277 603
rect 2282 543 2285 623
rect 2290 613 2293 643
rect 2250 413 2253 516
rect 2258 496 2261 526
rect 2274 523 2277 536
rect 2290 533 2293 606
rect 2298 573 2301 606
rect 2306 583 2309 616
rect 2258 493 2277 496
rect 2250 303 2253 316
rect 2258 223 2261 486
rect 2274 466 2277 493
rect 2282 473 2285 526
rect 2298 466 2301 526
rect 2274 463 2301 466
rect 2266 413 2269 446
rect 2274 403 2277 463
rect 2306 446 2309 546
rect 2302 443 2309 446
rect 2290 413 2293 436
rect 2302 386 2305 443
rect 2302 383 2309 386
rect 2266 216 2269 326
rect 2290 323 2293 346
rect 2298 313 2301 366
rect 2274 233 2277 306
rect 2306 223 2309 383
rect 2314 333 2317 1653
rect 2322 1613 2325 1706
rect 2330 1656 2333 1736
rect 2338 1693 2341 1813
rect 2346 1803 2357 1806
rect 2362 1793 2365 1806
rect 2354 1733 2357 1746
rect 2346 1723 2357 1726
rect 2362 1723 2365 1736
rect 2330 1653 2341 1656
rect 2346 1616 2349 1723
rect 2354 1663 2357 1716
rect 2370 1713 2373 1896
rect 2378 1873 2381 1926
rect 2394 1896 2397 1933
rect 2402 1903 2405 1963
rect 2410 1896 2413 1926
rect 2394 1893 2413 1896
rect 2418 1893 2421 1926
rect 2426 1906 2429 2233
rect 2450 2223 2453 2246
rect 2434 2193 2437 2216
rect 2458 2176 2461 2216
rect 2434 2173 2461 2176
rect 2434 2153 2437 2173
rect 2434 2133 2445 2136
rect 2434 1946 2437 2126
rect 2450 2063 2453 2136
rect 2442 2003 2445 2026
rect 2458 2013 2461 2166
rect 2466 2133 2469 2316
rect 2498 2296 2501 2343
rect 2514 2313 2517 2326
rect 2490 2293 2501 2296
rect 2474 2123 2477 2256
rect 2482 2193 2485 2206
rect 2482 2133 2485 2146
rect 2474 2043 2477 2076
rect 2466 2033 2477 2036
rect 2466 2003 2469 2033
rect 2482 2013 2485 2096
rect 2442 1993 2461 1996
rect 2434 1943 2445 1946
rect 2434 1923 2437 1936
rect 2426 1903 2433 1906
rect 2378 1823 2389 1826
rect 2386 1793 2389 1816
rect 2394 1723 2397 1836
rect 2402 1806 2405 1846
rect 2402 1803 2413 1806
rect 2418 1803 2421 1846
rect 2430 1836 2433 1903
rect 2442 1863 2445 1943
rect 2450 1923 2453 1936
rect 2458 1933 2461 1956
rect 2466 1906 2469 1996
rect 2474 1933 2477 1966
rect 2458 1903 2469 1906
rect 2474 1913 2485 1916
rect 2458 1873 2461 1903
rect 2474 1896 2477 1913
rect 2466 1893 2477 1896
rect 2466 1853 2469 1893
rect 2490 1886 2493 2293
rect 2514 2226 2517 2306
rect 2514 2223 2525 2226
rect 2498 2153 2501 2196
rect 2506 2146 2509 2206
rect 2514 2193 2517 2206
rect 2522 2193 2525 2223
rect 2498 2143 2517 2146
rect 2474 1883 2493 1886
rect 2474 1846 2477 1883
rect 2498 1876 2501 2136
rect 2514 2113 2517 2126
rect 2522 2093 2525 2136
rect 2506 2003 2509 2046
rect 2530 2026 2533 2356
rect 2538 2213 2541 2373
rect 2546 2363 2549 2416
rect 2562 2326 2565 2346
rect 2546 2293 2549 2326
rect 2558 2323 2565 2326
rect 2558 2246 2561 2323
rect 2570 2286 2573 2336
rect 2578 2303 2581 2416
rect 2586 2413 2597 2416
rect 2602 2413 2613 2416
rect 2586 2383 2589 2406
rect 2610 2403 2613 2413
rect 2618 2383 2621 2426
rect 2594 2333 2597 2346
rect 2570 2283 2597 2286
rect 2558 2243 2565 2246
rect 2546 2203 2549 2216
rect 2562 2203 2565 2243
rect 2538 2083 2541 2126
rect 2546 2076 2549 2176
rect 2562 2163 2573 2166
rect 2514 2023 2533 2026
rect 2538 2073 2549 2076
rect 2514 2013 2525 2016
rect 2514 1996 2517 2013
rect 2538 2006 2541 2073
rect 2546 2013 2549 2056
rect 2522 2003 2541 2006
rect 2554 2003 2557 2136
rect 2562 2083 2565 2136
rect 2570 2133 2573 2163
rect 2570 2113 2573 2126
rect 2578 2106 2581 2196
rect 2570 2103 2581 2106
rect 2514 1993 2533 1996
rect 2514 1983 2525 1986
rect 2506 1923 2509 1966
rect 2514 1883 2517 1916
rect 2426 1833 2433 1836
rect 2466 1843 2477 1846
rect 2386 1663 2389 1716
rect 2338 1613 2349 1616
rect 2322 1533 2325 1586
rect 2330 1553 2333 1606
rect 2330 1533 2333 1546
rect 2338 1526 2341 1613
rect 2330 1523 2341 1526
rect 2322 1493 2325 1516
rect 2330 1503 2333 1523
rect 2346 1473 2349 1606
rect 2354 1576 2357 1646
rect 2362 1583 2365 1656
rect 2394 1616 2397 1636
rect 2370 1603 2373 1616
rect 2378 1613 2397 1616
rect 2370 1586 2373 1596
rect 2394 1586 2397 1606
rect 2402 1593 2405 1736
rect 2410 1723 2413 1803
rect 2426 1756 2429 1833
rect 2442 1823 2453 1826
rect 2434 1813 2445 1816
rect 2426 1753 2433 1756
rect 2410 1596 2413 1626
rect 2418 1603 2421 1746
rect 2430 1626 2433 1753
rect 2442 1743 2445 1813
rect 2450 1793 2453 1823
rect 2458 1813 2461 1826
rect 2466 1813 2469 1843
rect 2458 1766 2461 1806
rect 2482 1773 2485 1876
rect 2494 1873 2501 1876
rect 2494 1806 2497 1873
rect 2490 1803 2497 1806
rect 2450 1763 2461 1766
rect 2450 1743 2461 1746
rect 2442 1703 2445 1736
rect 2450 1733 2453 1743
rect 2458 1706 2461 1726
rect 2458 1703 2465 1706
rect 2426 1623 2433 1626
rect 2410 1593 2421 1596
rect 2370 1583 2397 1586
rect 2354 1573 2365 1576
rect 2322 1083 2325 1416
rect 2338 1403 2341 1416
rect 2330 1323 2333 1336
rect 2346 1333 2349 1426
rect 2354 1293 2357 1546
rect 2362 1523 2365 1573
rect 2362 1493 2365 1516
rect 2362 1423 2365 1436
rect 2362 1386 2365 1406
rect 2370 1403 2373 1416
rect 2378 1403 2381 1566
rect 2394 1386 2397 1536
rect 2418 1526 2421 1593
rect 2426 1536 2429 1623
rect 2434 1546 2437 1606
rect 2450 1553 2453 1686
rect 2462 1626 2465 1703
rect 2474 1643 2477 1756
rect 2458 1623 2465 1626
rect 2458 1563 2461 1623
rect 2474 1606 2477 1626
rect 2482 1613 2485 1766
rect 2490 1733 2493 1803
rect 2498 1656 2501 1786
rect 2506 1726 2509 1806
rect 2514 1773 2517 1826
rect 2514 1733 2517 1766
rect 2506 1723 2517 1726
rect 2522 1723 2525 1983
rect 2530 1933 2533 1993
rect 2530 1903 2533 1926
rect 2498 1653 2509 1656
rect 2490 1613 2493 1636
rect 2466 1546 2469 1606
rect 2474 1603 2493 1606
rect 2506 1603 2509 1653
rect 2514 1603 2517 1723
rect 2530 1683 2533 1886
rect 2538 1873 2541 2003
rect 2546 1953 2549 1996
rect 2562 1983 2565 2016
rect 2546 1933 2557 1936
rect 2538 1833 2541 1856
rect 2546 1826 2549 1916
rect 2562 1856 2565 1926
rect 2570 1923 2573 2103
rect 2578 2043 2581 2076
rect 2578 2023 2581 2036
rect 2562 1853 2573 1856
rect 2538 1823 2549 1826
rect 2554 1823 2557 1836
rect 2538 1806 2541 1823
rect 2546 1813 2557 1816
rect 2538 1803 2545 1806
rect 2542 1736 2545 1803
rect 2554 1783 2557 1813
rect 2542 1733 2549 1736
rect 2538 1676 2541 1716
rect 2522 1673 2541 1676
rect 2522 1606 2525 1673
rect 2530 1613 2533 1666
rect 2522 1603 2529 1606
rect 2490 1546 2493 1603
rect 2434 1543 2453 1546
rect 2426 1533 2437 1536
rect 2410 1503 2413 1526
rect 2418 1523 2429 1526
rect 2434 1516 2437 1533
rect 2426 1513 2437 1516
rect 2410 1393 2413 1426
rect 2362 1383 2373 1386
rect 2370 1286 2373 1383
rect 2386 1383 2397 1386
rect 2386 1366 2389 1383
rect 2362 1283 2373 1286
rect 2382 1363 2389 1366
rect 2362 1266 2365 1283
rect 2358 1263 2365 1266
rect 2330 1216 2333 1226
rect 2330 1213 2341 1216
rect 2330 1063 2333 1206
rect 2338 1106 2341 1213
rect 2358 1206 2361 1263
rect 2382 1246 2385 1363
rect 2382 1243 2389 1246
rect 2354 1203 2361 1206
rect 2354 1173 2357 1203
rect 2370 1186 2373 1236
rect 2386 1223 2389 1243
rect 2366 1183 2373 1186
rect 2346 1123 2349 1136
rect 2354 1133 2357 1156
rect 2338 1103 2345 1106
rect 2342 1036 2345 1103
rect 2338 1033 2345 1036
rect 2322 983 2325 996
rect 2330 963 2333 1016
rect 2322 843 2325 946
rect 2338 943 2341 1033
rect 2354 936 2357 1126
rect 2366 956 2369 1183
rect 2378 1143 2381 1196
rect 2366 953 2373 956
rect 2354 933 2365 936
rect 2338 853 2341 926
rect 2322 816 2325 826
rect 2322 813 2333 816
rect 2322 793 2325 806
rect 2338 803 2341 846
rect 2346 786 2349 816
rect 2354 803 2357 926
rect 2362 823 2365 933
rect 2362 793 2365 816
rect 2342 783 2349 786
rect 2330 736 2333 776
rect 2322 733 2333 736
rect 2342 726 2345 783
rect 2370 766 2373 953
rect 2378 923 2381 1136
rect 2386 1003 2389 1206
rect 2394 1166 2397 1376
rect 2402 1313 2405 1336
rect 2418 1333 2421 1346
rect 2418 1303 2421 1326
rect 2402 1213 2405 1226
rect 2410 1213 2413 1236
rect 2410 1203 2421 1206
rect 2418 1183 2421 1203
rect 2394 1163 2405 1166
rect 2402 1076 2405 1163
rect 2426 1146 2429 1513
rect 2442 1493 2445 1526
rect 2442 1373 2445 1416
rect 2450 1346 2453 1543
rect 2458 1543 2469 1546
rect 2458 1506 2461 1543
rect 2466 1513 2469 1536
rect 2458 1503 2465 1506
rect 2462 1426 2465 1503
rect 2462 1423 2469 1426
rect 2458 1383 2461 1396
rect 2442 1343 2453 1346
rect 2434 1323 2437 1336
rect 2442 1323 2445 1343
rect 2434 1213 2437 1226
rect 2442 1203 2445 1286
rect 2450 1183 2453 1336
rect 2458 1313 2461 1326
rect 2466 1303 2469 1423
rect 2394 1073 2405 1076
rect 2418 1143 2429 1146
rect 2394 1003 2397 1073
rect 2394 933 2397 996
rect 2402 993 2405 1056
rect 2418 1026 2421 1143
rect 2418 1023 2429 1026
rect 2410 1003 2421 1006
rect 2418 953 2421 996
rect 2378 803 2381 856
rect 2370 763 2381 766
rect 2354 733 2357 756
rect 2370 743 2373 756
rect 2342 723 2349 726
rect 2322 626 2325 646
rect 2346 636 2349 723
rect 2342 633 2349 636
rect 2322 623 2333 626
rect 2330 556 2333 623
rect 2322 553 2333 556
rect 2342 556 2345 633
rect 2354 593 2357 626
rect 2342 553 2349 556
rect 2322 413 2325 553
rect 2330 386 2333 526
rect 2338 473 2341 536
rect 2322 383 2333 386
rect 2322 333 2325 383
rect 2314 223 2325 226
rect 2266 213 2317 216
rect 2234 203 2253 206
rect 2194 173 2205 176
rect 2202 126 2205 173
rect 2250 143 2253 203
rect 2266 136 2269 213
rect 2226 133 2245 136
rect 2194 123 2205 126
rect 2194 103 2197 123
rect 2242 53 2245 133
rect 2250 133 2269 136
rect 2298 133 2301 206
rect 2322 193 2325 223
rect 2250 123 2253 133
rect 2314 66 2317 126
rect 2306 63 2317 66
rect 2322 63 2325 136
rect 2330 103 2333 376
rect 2346 336 2349 553
rect 2354 343 2357 546
rect 2362 386 2365 726
rect 2370 713 2373 736
rect 2370 553 2373 616
rect 2378 536 2381 763
rect 2386 623 2389 896
rect 2402 866 2405 926
rect 2410 893 2413 936
rect 2418 933 2421 946
rect 2394 863 2405 866
rect 2394 763 2397 796
rect 2410 773 2413 866
rect 2418 853 2421 926
rect 2426 836 2429 1023
rect 2434 933 2437 1136
rect 2442 1096 2445 1126
rect 2450 1123 2453 1136
rect 2458 1123 2461 1296
rect 2474 1216 2477 1546
rect 2490 1543 2501 1546
rect 2482 1503 2485 1526
rect 2498 1523 2501 1543
rect 2498 1416 2501 1436
rect 2482 1413 2501 1416
rect 2482 1306 2485 1413
rect 2498 1346 2501 1406
rect 2490 1343 2501 1346
rect 2490 1323 2493 1343
rect 2482 1303 2493 1306
rect 2490 1236 2493 1303
rect 2466 1213 2477 1216
rect 2482 1233 2493 1236
rect 2466 1173 2469 1213
rect 2482 1156 2485 1233
rect 2498 1196 2501 1216
rect 2474 1153 2485 1156
rect 2494 1193 2501 1196
rect 2474 1106 2477 1153
rect 2494 1116 2497 1193
rect 2506 1123 2509 1596
rect 2526 1546 2529 1603
rect 2514 1533 2517 1546
rect 2526 1543 2533 1546
rect 2514 1413 2517 1516
rect 2522 1453 2525 1526
rect 2530 1373 2533 1543
rect 2538 1533 2541 1626
rect 2538 1503 2541 1526
rect 2546 1486 2549 1733
rect 2554 1706 2557 1736
rect 2562 1723 2565 1826
rect 2570 1823 2573 1853
rect 2578 1823 2581 2016
rect 2586 1996 2589 2276
rect 2594 2193 2597 2283
rect 2610 2213 2613 2296
rect 2626 2256 2629 2396
rect 2642 2353 2645 2443
rect 2666 2386 2669 2443
rect 2662 2383 2669 2386
rect 2642 2323 2645 2346
rect 2626 2253 2633 2256
rect 2630 2196 2633 2253
rect 2642 2203 2645 2216
rect 2650 2203 2653 2276
rect 2662 2256 2665 2383
rect 2674 2283 2677 2516
rect 2682 2293 2685 2553
rect 2690 2393 2693 2416
rect 2714 2386 2717 2526
rect 2730 2513 2733 2563
rect 2738 2533 2741 2606
rect 2746 2533 2749 2606
rect 2754 2506 2757 2526
rect 2738 2503 2757 2506
rect 2738 2436 2741 2503
rect 2730 2433 2741 2436
rect 2730 2396 2733 2433
rect 2762 2423 2765 2616
rect 2778 2613 2781 2716
rect 2810 2656 2813 2736
rect 2818 2713 2821 2726
rect 2834 2703 2837 2716
rect 2842 2656 2845 2816
rect 2850 2776 2853 2963
rect 2882 2923 2885 2936
rect 2898 2933 2901 3196
rect 2930 3156 2933 3216
rect 2922 3153 2933 3156
rect 2922 3013 2925 3153
rect 2946 3123 2949 3216
rect 2970 3183 2973 3206
rect 3018 3176 3021 3216
rect 3074 3213 3077 3253
rect 3114 3213 3117 3253
rect 3290 3253 3333 3256
rect 3090 3193 3093 3206
rect 3018 3173 3029 3176
rect 2986 3133 2989 3146
rect 3026 3133 3029 3173
rect 2938 2923 2941 3016
rect 2946 3013 2949 3026
rect 2954 2996 2957 3006
rect 2978 3003 2981 3126
rect 3034 3106 3037 3126
rect 3042 3116 3045 3146
rect 3058 3133 3061 3156
rect 3050 3123 3061 3126
rect 3066 3116 3069 3126
rect 3074 3123 3085 3126
rect 3042 3113 3069 3116
rect 3026 3103 3037 3106
rect 3026 3046 3029 3103
rect 3082 3076 3085 3116
rect 3050 3073 3085 3076
rect 3026 3043 3037 3046
rect 3002 3023 3029 3026
rect 3034 3023 3037 3043
rect 3002 2996 3005 3006
rect 3010 3003 3013 3016
rect 2954 2993 3005 2996
rect 2970 2926 2973 2986
rect 3018 2976 3021 3016
rect 3026 3006 3029 3023
rect 3026 3003 3037 3006
rect 2994 2973 3021 2976
rect 2994 2926 2997 2973
rect 3042 2926 3045 3016
rect 2970 2923 2997 2926
rect 3010 2923 3045 2926
rect 2986 2856 2989 2916
rect 2994 2903 2997 2923
rect 3050 2916 3053 3073
rect 3106 3033 3109 3136
rect 3122 3133 3133 3136
rect 3138 3073 3141 3146
rect 3114 3043 3157 3046
rect 3082 3023 3109 3026
rect 3114 3023 3117 3043
rect 3082 3013 3085 3023
rect 3106 3016 3109 3023
rect 3058 2983 3061 3006
rect 3074 3003 3085 3006
rect 3074 2996 3077 3003
rect 3066 2993 3077 2996
rect 3066 2933 3069 2993
rect 3082 2926 3085 2996
rect 3098 2993 3101 3016
rect 3106 3013 3117 3016
rect 3074 2923 3085 2926
rect 3002 2913 3029 2916
rect 3042 2913 3053 2916
rect 2978 2853 2989 2856
rect 2850 2773 2857 2776
rect 2810 2653 2845 2656
rect 2818 2613 2821 2626
rect 2770 2523 2773 2606
rect 2778 2533 2781 2606
rect 2786 2576 2789 2606
rect 2834 2603 2837 2636
rect 2786 2573 2793 2576
rect 2790 2526 2793 2573
rect 2786 2523 2793 2526
rect 2786 2426 2789 2523
rect 2810 2513 2813 2536
rect 2842 2533 2845 2653
rect 2854 2636 2857 2773
rect 2850 2633 2857 2636
rect 2850 2613 2853 2633
rect 2866 2576 2869 2806
rect 2890 2756 2893 2816
rect 2946 2813 2949 2826
rect 2978 2803 2981 2853
rect 2994 2816 2997 2826
rect 3002 2823 3005 2913
rect 3026 2903 3037 2906
rect 2986 2813 3005 2816
rect 3026 2776 3029 2836
rect 3050 2803 3053 2876
rect 3026 2773 3037 2776
rect 2882 2753 2893 2756
rect 2882 2706 2885 2753
rect 2898 2743 2941 2746
rect 2898 2716 2901 2726
rect 2898 2713 2917 2716
rect 2882 2703 2893 2706
rect 2890 2643 2893 2703
rect 2874 2613 2877 2626
rect 2882 2593 2885 2616
rect 2850 2573 2869 2576
rect 2850 2526 2853 2573
rect 2890 2543 2893 2606
rect 2842 2523 2853 2526
rect 2858 2523 2861 2536
rect 2786 2423 2813 2426
rect 2738 2406 2741 2416
rect 2746 2413 2781 2416
rect 2738 2403 2757 2406
rect 2730 2393 2749 2396
rect 2706 2383 2733 2386
rect 2706 2333 2709 2383
rect 2730 2333 2733 2346
rect 2738 2333 2741 2356
rect 2690 2273 2693 2326
rect 2714 2323 2733 2326
rect 2746 2316 2749 2393
rect 2754 2376 2757 2403
rect 2762 2393 2765 2406
rect 2754 2373 2761 2376
rect 2730 2313 2749 2316
rect 2758 2306 2761 2373
rect 2770 2363 2773 2406
rect 2754 2303 2761 2306
rect 2662 2253 2669 2256
rect 2666 2233 2669 2253
rect 2682 2213 2685 2266
rect 2738 2226 2741 2256
rect 2698 2213 2701 2226
rect 2706 2223 2741 2226
rect 2626 2193 2633 2196
rect 2626 2173 2629 2193
rect 2594 2093 2597 2116
rect 2594 2013 2597 2076
rect 2586 1993 2593 1996
rect 2590 1926 2593 1993
rect 2590 1923 2597 1926
rect 2586 1883 2589 1916
rect 2594 1873 2597 1923
rect 2602 1836 2605 2136
rect 2610 2123 2613 2166
rect 2610 2043 2613 2056
rect 2618 2036 2621 2136
rect 2634 2123 2637 2136
rect 2642 2133 2645 2146
rect 2658 2126 2661 2136
rect 2642 2113 2645 2126
rect 2650 2123 2661 2126
rect 2650 2053 2653 2123
rect 2658 2036 2661 2116
rect 2578 1783 2581 1816
rect 2586 1803 2589 1836
rect 2594 1833 2605 1836
rect 2610 2033 2621 2036
rect 2626 2033 2661 2036
rect 2570 1733 2573 1756
rect 2578 1723 2589 1726
rect 2554 1703 2561 1706
rect 2558 1636 2561 1703
rect 2542 1483 2549 1486
rect 2554 1633 2561 1636
rect 2554 1483 2557 1633
rect 2562 1573 2565 1616
rect 2542 1416 2545 1483
rect 2542 1413 2549 1416
rect 2514 1306 2517 1336
rect 2530 1333 2533 1346
rect 2538 1326 2541 1396
rect 2522 1323 2541 1326
rect 2546 1306 2549 1413
rect 2514 1303 2525 1306
rect 2522 1236 2525 1303
rect 2538 1303 2549 1306
rect 2538 1246 2541 1303
rect 2538 1243 2549 1246
rect 2514 1233 2525 1236
rect 2514 1213 2517 1233
rect 2522 1213 2533 1216
rect 2514 1133 2517 1196
rect 2494 1113 2501 1116
rect 2474 1103 2485 1106
rect 2442 1093 2461 1096
rect 2466 1016 2469 1036
rect 2450 1013 2469 1016
rect 2450 986 2453 1013
rect 2442 983 2453 986
rect 2434 903 2437 926
rect 2434 853 2437 896
rect 2422 833 2429 836
rect 2394 733 2397 746
rect 2422 736 2425 833
rect 2442 813 2445 983
rect 2434 753 2437 806
rect 2450 746 2453 936
rect 2434 743 2453 746
rect 2458 736 2461 966
rect 2482 963 2485 1103
rect 2498 1026 2501 1113
rect 2522 1073 2525 1213
rect 2530 1183 2533 1206
rect 2538 1203 2541 1226
rect 2530 1133 2541 1136
rect 2530 1123 2541 1126
rect 2546 1106 2549 1243
rect 2554 1213 2557 1446
rect 2562 1423 2565 1536
rect 2538 1103 2549 1106
rect 2538 1036 2541 1103
rect 2538 1033 2549 1036
rect 2494 1023 2501 1026
rect 2494 956 2497 1023
rect 2546 1016 2549 1033
rect 2506 1013 2533 1016
rect 2522 976 2525 1006
rect 2530 1003 2533 1013
rect 2538 1013 2549 1016
rect 2506 973 2525 976
rect 2494 953 2501 956
rect 2466 933 2469 946
rect 2474 933 2493 936
rect 2466 833 2469 866
rect 2394 703 2397 726
rect 2402 723 2405 736
rect 2422 733 2429 736
rect 2394 613 2397 646
rect 2370 533 2381 536
rect 2370 496 2373 533
rect 2378 513 2381 526
rect 2394 503 2397 576
rect 2370 493 2381 496
rect 2378 426 2381 493
rect 2402 446 2405 536
rect 2410 523 2413 666
rect 2418 583 2421 606
rect 2426 526 2429 733
rect 2450 733 2461 736
rect 2466 733 2469 826
rect 2434 533 2437 626
rect 2442 583 2445 616
rect 2426 523 2437 526
rect 2402 443 2421 446
rect 2370 423 2381 426
rect 2370 403 2373 423
rect 2362 383 2373 386
rect 2346 333 2357 336
rect 2338 213 2341 226
rect 2346 223 2349 326
rect 2354 316 2357 333
rect 2354 313 2361 316
rect 2358 256 2361 313
rect 2354 253 2361 256
rect 2354 203 2357 253
rect 2370 236 2373 383
rect 2386 303 2389 346
rect 2394 313 2397 416
rect 2410 413 2413 436
rect 2402 286 2405 406
rect 2410 303 2413 316
rect 2418 313 2421 443
rect 2426 423 2429 466
rect 2434 413 2437 523
rect 2426 393 2437 396
rect 2426 323 2429 393
rect 2442 386 2445 486
rect 2434 383 2445 386
rect 2402 283 2413 286
rect 2362 233 2373 236
rect 2362 183 2365 233
rect 2386 223 2389 236
rect 2394 223 2397 266
rect 2410 216 2413 283
rect 2378 183 2381 216
rect 2402 213 2413 216
rect 2346 113 2349 136
rect 2378 133 2381 166
rect 2402 123 2405 213
rect 2434 203 2437 383
rect 2450 306 2453 733
rect 2466 706 2469 726
rect 2458 703 2469 706
rect 2474 686 2477 933
rect 2490 853 2493 916
rect 2498 836 2501 953
rect 2506 943 2509 973
rect 2506 923 2509 936
rect 2506 863 2509 916
rect 2494 833 2501 836
rect 2470 683 2477 686
rect 2470 626 2473 683
rect 2470 623 2477 626
rect 2458 533 2461 606
rect 2458 443 2461 526
rect 2466 376 2469 606
rect 2474 466 2477 623
rect 2482 586 2485 816
rect 2494 786 2497 833
rect 2506 793 2509 836
rect 2514 803 2517 966
rect 2538 963 2541 1013
rect 2546 993 2549 1006
rect 2522 933 2533 936
rect 2538 933 2541 946
rect 2494 783 2501 786
rect 2498 736 2501 783
rect 2490 733 2501 736
rect 2514 726 2517 736
rect 2506 723 2517 726
rect 2490 603 2493 626
rect 2498 623 2501 656
rect 2482 583 2489 586
rect 2486 516 2489 583
rect 2498 533 2501 586
rect 2506 543 2509 723
rect 2522 713 2525 906
rect 2546 843 2549 926
rect 2554 863 2557 1206
rect 2562 1173 2565 1266
rect 2562 1123 2565 1136
rect 2562 923 2565 1076
rect 2570 1013 2573 1716
rect 2578 1463 2581 1696
rect 2594 1663 2597 1833
rect 2586 1546 2589 1596
rect 2594 1553 2597 1616
rect 2602 1613 2605 1826
rect 2610 1823 2613 2033
rect 2626 2006 2629 2033
rect 2618 2003 2629 2006
rect 2618 1916 2621 2003
rect 2626 1923 2629 1966
rect 2634 1946 2637 2006
rect 2642 1983 2645 2016
rect 2658 2006 2661 2026
rect 2666 2013 2669 2166
rect 2634 1943 2645 1946
rect 2650 1943 2653 2006
rect 2658 2003 2669 2006
rect 2666 1943 2669 2003
rect 2618 1913 2629 1916
rect 2642 1913 2645 1926
rect 2618 1883 2621 1906
rect 2610 1693 2613 1736
rect 2618 1713 2621 1876
rect 2626 1833 2629 1913
rect 2650 1906 2653 1936
rect 2634 1903 2653 1906
rect 2658 1933 2669 1936
rect 2658 1896 2661 1933
rect 2650 1893 2661 1896
rect 2650 1833 2653 1893
rect 2634 1803 2637 1826
rect 2658 1823 2661 1856
rect 2666 1803 2669 1926
rect 2674 1813 2677 2176
rect 2698 2156 2701 2206
rect 2706 2203 2709 2223
rect 2714 2203 2717 2216
rect 2722 2163 2725 2223
rect 2730 2156 2733 2216
rect 2698 2153 2733 2156
rect 2682 2106 2685 2126
rect 2682 2103 2689 2106
rect 2686 2036 2689 2103
rect 2698 2083 2701 2116
rect 2706 2093 2709 2126
rect 2682 2033 2689 2036
rect 2682 2016 2685 2033
rect 2682 2013 2693 2016
rect 2682 1933 2685 1976
rect 2690 1943 2693 1996
rect 2698 1936 2701 2046
rect 2706 1943 2709 2026
rect 2698 1933 2709 1936
rect 2682 1923 2701 1926
rect 2682 1806 2685 1826
rect 2674 1803 2685 1806
rect 2626 1726 2629 1756
rect 2634 1733 2653 1736
rect 2658 1733 2661 1746
rect 2626 1723 2637 1726
rect 2610 1583 2613 1606
rect 2618 1603 2621 1616
rect 2626 1596 2629 1696
rect 2634 1613 2637 1723
rect 2618 1593 2629 1596
rect 2634 1593 2637 1606
rect 2586 1543 2597 1546
rect 2586 1523 2589 1536
rect 2594 1456 2597 1543
rect 2578 1453 2597 1456
rect 2578 1393 2581 1453
rect 2602 1443 2605 1526
rect 2594 1413 2597 1436
rect 2602 1413 2605 1426
rect 2610 1376 2613 1466
rect 2594 1373 2613 1376
rect 2586 1223 2589 1356
rect 2594 1223 2597 1373
rect 2602 1293 2605 1336
rect 2610 1273 2613 1336
rect 2618 1256 2621 1593
rect 2642 1583 2645 1726
rect 2650 1603 2653 1733
rect 2658 1713 2661 1726
rect 2666 1716 2669 1776
rect 2674 1743 2677 1803
rect 2682 1736 2685 1766
rect 2690 1743 2693 1886
rect 2698 1873 2701 1923
rect 2706 1883 2709 1933
rect 2714 1906 2717 2136
rect 2722 2043 2725 2136
rect 2722 1923 2725 2026
rect 2730 2013 2733 2106
rect 2714 1903 2721 1906
rect 2698 1833 2701 1846
rect 2682 1733 2693 1736
rect 2690 1723 2693 1733
rect 2698 1716 2701 1826
rect 2706 1723 2709 1866
rect 2718 1826 2721 1903
rect 2730 1853 2733 2006
rect 2738 1836 2741 2216
rect 2746 2133 2749 2226
rect 2754 2203 2757 2303
rect 2770 2213 2773 2346
rect 2778 2323 2781 2413
rect 2786 2393 2789 2406
rect 2794 2333 2797 2416
rect 2810 2363 2813 2423
rect 2810 2333 2813 2356
rect 2786 2313 2805 2316
rect 2786 2213 2789 2246
rect 2802 2213 2805 2313
rect 2818 2246 2821 2326
rect 2826 2263 2829 2416
rect 2842 2403 2845 2523
rect 2882 2486 2885 2506
rect 2878 2483 2885 2486
rect 2866 2353 2869 2416
rect 2878 2386 2881 2483
rect 2878 2383 2885 2386
rect 2874 2346 2877 2366
rect 2834 2343 2877 2346
rect 2882 2343 2885 2383
rect 2834 2333 2837 2343
rect 2842 2293 2845 2336
rect 2810 2243 2821 2246
rect 2850 2243 2853 2336
rect 2858 2333 2869 2336
rect 2874 2333 2877 2343
rect 2746 2013 2749 2086
rect 2754 2006 2757 2196
rect 2762 2113 2765 2176
rect 2770 2076 2773 2166
rect 2770 2073 2789 2076
rect 2762 2013 2765 2056
rect 2746 2003 2757 2006
rect 2746 1943 2749 2003
rect 2762 1963 2765 2006
rect 2770 1956 2773 2066
rect 2786 2063 2789 2073
rect 2778 1983 2781 2016
rect 2786 2003 2789 2036
rect 2770 1953 2789 1956
rect 2746 1933 2757 1936
rect 2746 1896 2749 1933
rect 2754 1913 2757 1926
rect 2762 1903 2765 1936
rect 2770 1923 2773 1946
rect 2786 1933 2789 1953
rect 2778 1923 2789 1926
rect 2746 1893 2753 1896
rect 2714 1823 2721 1826
rect 2730 1833 2741 1836
rect 2666 1713 2677 1716
rect 2690 1713 2701 1716
rect 2658 1596 2661 1706
rect 2674 1636 2677 1713
rect 2650 1593 2661 1596
rect 2666 1633 2677 1636
rect 2666 1596 2669 1633
rect 2690 1623 2701 1626
rect 2690 1603 2693 1623
rect 2666 1593 2677 1596
rect 2642 1506 2645 1546
rect 2650 1523 2653 1593
rect 2642 1503 2649 1506
rect 2614 1253 2621 1256
rect 2578 1203 2581 1216
rect 2570 916 2573 946
rect 2578 933 2581 1176
rect 2586 1153 2589 1216
rect 2586 1093 2589 1126
rect 2594 1103 2597 1216
rect 2602 1133 2605 1206
rect 2614 1146 2617 1253
rect 2626 1213 2629 1456
rect 2634 1223 2637 1496
rect 2646 1426 2649 1503
rect 2642 1423 2649 1426
rect 2634 1166 2637 1216
rect 2626 1163 2637 1166
rect 2614 1143 2621 1146
rect 2602 1076 2605 1126
rect 2586 1073 2605 1076
rect 2562 913 2573 916
rect 2530 823 2557 826
rect 2530 693 2533 726
rect 2514 533 2517 616
rect 2538 613 2541 796
rect 2554 793 2557 823
rect 2562 723 2565 913
rect 2578 903 2581 926
rect 2586 896 2589 1073
rect 2594 1003 2597 1016
rect 2602 976 2605 1066
rect 2610 1003 2613 1126
rect 2618 1073 2621 1143
rect 2626 1063 2629 1163
rect 2634 1133 2637 1156
rect 2642 1066 2645 1423
rect 2650 1393 2653 1406
rect 2650 1113 2653 1386
rect 2658 1323 2661 1586
rect 2666 1533 2669 1586
rect 2658 1203 2661 1256
rect 2658 1143 2661 1156
rect 2658 1083 2661 1136
rect 2642 1063 2649 1066
rect 2626 983 2629 1006
rect 2602 973 2629 976
rect 2570 893 2589 896
rect 2570 733 2573 893
rect 2594 886 2597 936
rect 2586 883 2597 886
rect 2578 753 2581 876
rect 2586 803 2589 883
rect 2594 813 2597 866
rect 2594 763 2597 806
rect 2602 796 2605 966
rect 2610 813 2613 946
rect 2618 916 2621 936
rect 2626 926 2629 973
rect 2634 956 2637 1056
rect 2646 1016 2649 1063
rect 2642 1013 2649 1016
rect 2642 963 2645 1013
rect 2634 953 2645 956
rect 2642 933 2645 953
rect 2650 926 2653 996
rect 2658 943 2661 1016
rect 2666 936 2669 1516
rect 2674 1453 2677 1593
rect 2674 1416 2677 1436
rect 2682 1426 2685 1576
rect 2690 1523 2693 1586
rect 2682 1423 2693 1426
rect 2674 1413 2693 1416
rect 2674 1333 2677 1376
rect 2682 1323 2685 1406
rect 2674 1083 2677 1316
rect 2682 1173 2685 1216
rect 2690 1213 2693 1413
rect 2698 1343 2701 1616
rect 2698 1213 2701 1256
rect 2706 1206 2709 1716
rect 2714 1583 2717 1823
rect 2722 1616 2725 1806
rect 2730 1776 2733 1833
rect 2738 1783 2741 1826
rect 2750 1796 2753 1893
rect 2778 1866 2781 1923
rect 2770 1863 2781 1866
rect 2762 1796 2765 1826
rect 2770 1823 2773 1863
rect 2778 1813 2781 1846
rect 2786 1836 2789 1916
rect 2794 1846 2797 2116
rect 2802 1873 2805 2206
rect 2810 2203 2813 2216
rect 2818 2173 2821 2243
rect 2834 2213 2837 2226
rect 2842 2206 2845 2236
rect 2826 2193 2829 2206
rect 2838 2203 2845 2206
rect 2838 2146 2841 2203
rect 2810 2096 2813 2146
rect 2818 2143 2829 2146
rect 2834 2143 2841 2146
rect 2850 2143 2853 2156
rect 2858 2146 2861 2333
rect 2866 2303 2869 2326
rect 2890 2253 2893 2526
rect 2898 2516 2901 2616
rect 2914 2613 2917 2713
rect 2922 2693 2925 2726
rect 2930 2656 2933 2736
rect 2938 2663 2941 2743
rect 2954 2713 2965 2716
rect 2930 2653 2973 2656
rect 2906 2553 2909 2606
rect 2922 2596 2925 2626
rect 2930 2603 2933 2653
rect 2914 2593 2925 2596
rect 2906 2523 2909 2536
rect 2914 2526 2917 2593
rect 2954 2586 2957 2646
rect 2962 2623 2965 2636
rect 2962 2593 2965 2606
rect 2970 2596 2973 2653
rect 2978 2623 2989 2626
rect 2970 2593 2981 2596
rect 2954 2583 2965 2586
rect 2922 2533 2933 2536
rect 2914 2523 2933 2526
rect 2898 2513 2933 2516
rect 2938 2503 2941 2536
rect 2962 2533 2965 2583
rect 2986 2556 2989 2616
rect 2994 2603 2997 2666
rect 3010 2643 3013 2716
rect 3018 2713 3021 2736
rect 3018 2613 3021 2696
rect 3034 2676 3037 2773
rect 3058 2753 3061 2916
rect 3074 2873 3077 2923
rect 3082 2903 3085 2916
rect 3090 2836 3093 2916
rect 3082 2833 3093 2836
rect 3066 2813 3069 2826
rect 3082 2823 3085 2833
rect 3098 2826 3101 2926
rect 3106 2903 3109 3006
rect 3114 2923 3117 3013
rect 3122 2963 3125 3036
rect 3130 3006 3133 3026
rect 3138 3013 3141 3036
rect 3130 3003 3141 3006
rect 3130 2993 3141 2996
rect 3138 2943 3141 2993
rect 3154 2976 3157 3043
rect 3170 2983 3173 3156
rect 3178 3133 3181 3216
rect 3202 3173 3205 3206
rect 3194 3133 3221 3136
rect 3250 3133 3253 3216
rect 3290 3213 3293 3253
rect 3330 3213 3333 3253
rect 3178 3123 3213 3126
rect 3210 3023 3213 3046
rect 3210 3003 3213 3016
rect 3218 2993 3221 3133
rect 3266 3126 3269 3136
rect 3290 3133 3293 3166
rect 3226 3086 3229 3126
rect 3266 3123 3293 3126
rect 3226 3083 3237 3086
rect 3226 3013 3229 3076
rect 3234 2986 3237 3083
rect 3242 3003 3245 3046
rect 3250 2996 3253 3006
rect 3226 2983 3237 2986
rect 3242 2993 3253 2996
rect 3154 2973 3173 2976
rect 3114 2913 3133 2916
rect 3090 2823 3101 2826
rect 3114 2823 3117 2913
rect 3138 2883 3141 2936
rect 3146 2933 3157 2936
rect 3154 2903 3157 2926
rect 3170 2923 3173 2973
rect 3202 2923 3205 2946
rect 3210 2933 3221 2936
rect 3226 2933 3229 2983
rect 3234 2933 3237 2946
rect 3242 2943 3245 2993
rect 3258 2966 3261 3076
rect 3274 3013 3277 3123
rect 3282 3113 3293 3116
rect 3298 3073 3301 3136
rect 3306 3036 3309 3206
rect 3314 3143 3317 3166
rect 3386 3153 3389 3216
rect 3314 3116 3317 3136
rect 3354 3123 3357 3136
rect 3314 3113 3325 3116
rect 3322 3066 3325 3113
rect 3250 2963 3261 2966
rect 3218 2913 3221 2926
rect 3242 2923 3245 2936
rect 3250 2926 3253 2963
rect 3266 2956 3269 3006
rect 3258 2953 3269 2956
rect 3258 2933 3261 2953
rect 3274 2946 3277 3006
rect 3282 3003 3285 3036
rect 3298 3033 3309 3036
rect 3314 3063 3325 3066
rect 3298 2986 3301 3033
rect 3314 3013 3317 3063
rect 3314 2986 3317 3006
rect 3354 3003 3357 3016
rect 3394 3013 3397 3076
rect 3298 2983 3317 2986
rect 3266 2943 3277 2946
rect 3298 2963 3341 2966
rect 3298 2933 3301 2963
rect 3250 2923 3261 2926
rect 3258 2903 3261 2923
rect 3282 2913 3285 2926
rect 3314 2893 3317 2936
rect 3338 2923 3341 2963
rect 3394 2923 3397 3006
rect 3090 2746 3093 2823
rect 3098 2813 3117 2816
rect 3194 2813 3197 2826
rect 3210 2813 3221 2816
rect 3178 2793 3181 2806
rect 3066 2733 3069 2746
rect 3090 2743 3101 2746
rect 3050 2693 3053 2726
rect 3098 2696 3101 2743
rect 3162 2733 3165 2746
rect 3194 2736 3197 2806
rect 3202 2793 3205 2806
rect 3218 2766 3221 2806
rect 3226 2803 3229 2836
rect 3234 2806 3237 2816
rect 3290 2813 3309 2816
rect 3314 2813 3333 2816
rect 3234 2803 3253 2806
rect 3274 2803 3293 2806
rect 3218 2763 3233 2766
rect 3194 2733 3201 2736
rect 3090 2693 3101 2696
rect 3034 2673 3045 2676
rect 3042 2616 3045 2673
rect 3090 2626 3093 2693
rect 3114 2686 3117 2726
rect 3146 2713 3149 2726
rect 3114 2683 3133 2686
rect 3130 2666 3133 2683
rect 3130 2663 3137 2666
rect 3026 2613 3045 2616
rect 3086 2623 3093 2626
rect 3106 2653 3125 2656
rect 2978 2553 2989 2556
rect 2946 2513 2965 2516
rect 2874 2203 2877 2216
rect 2858 2143 2877 2146
rect 2826 2123 2829 2136
rect 2810 2093 2821 2096
rect 2810 2023 2813 2086
rect 2794 1843 2805 1846
rect 2786 1833 2797 1836
rect 2786 1806 2789 1826
rect 2770 1803 2789 1806
rect 2750 1793 2773 1796
rect 2746 1783 2757 1786
rect 2730 1773 2749 1776
rect 2754 1773 2757 1783
rect 2730 1693 2733 1766
rect 2738 1733 2741 1746
rect 2730 1623 2733 1646
rect 2722 1613 2733 1616
rect 2714 1463 2717 1526
rect 2722 1433 2725 1596
rect 2730 1523 2733 1556
rect 2738 1493 2741 1726
rect 2746 1603 2749 1773
rect 2762 1723 2765 1793
rect 2754 1713 2765 1716
rect 2754 1696 2757 1713
rect 2754 1693 2761 1696
rect 2758 1626 2761 1693
rect 2754 1623 2761 1626
rect 2714 1413 2717 1426
rect 2738 1423 2741 1466
rect 2722 1413 2733 1416
rect 2714 1393 2717 1406
rect 2714 1333 2717 1346
rect 2698 1203 2709 1206
rect 2698 1156 2701 1203
rect 2690 1133 2693 1156
rect 2698 1153 2709 1156
rect 2682 1123 2693 1126
rect 2674 973 2677 1066
rect 2682 1013 2685 1123
rect 2682 943 2685 1006
rect 2626 923 2637 926
rect 2642 923 2653 926
rect 2642 916 2645 923
rect 2618 913 2645 916
rect 2658 906 2661 936
rect 2666 933 2685 936
rect 2602 793 2609 796
rect 2594 726 2597 736
rect 2586 723 2597 726
rect 2562 703 2565 716
rect 2522 543 2525 606
rect 2546 546 2549 616
rect 2554 603 2557 676
rect 2586 646 2589 723
rect 2594 703 2597 716
rect 2606 696 2609 793
rect 2618 723 2621 866
rect 2634 793 2637 906
rect 2650 903 2661 906
rect 2666 906 2669 926
rect 2666 903 2673 906
rect 2578 643 2589 646
rect 2602 693 2609 696
rect 2562 613 2565 636
rect 2530 543 2549 546
rect 2482 513 2489 516
rect 2482 493 2485 513
rect 2474 463 2485 466
rect 2474 413 2477 456
rect 2482 383 2485 463
rect 2498 456 2501 526
rect 2506 483 2509 526
rect 2530 456 2533 543
rect 2538 493 2541 526
rect 2546 513 2549 536
rect 2554 523 2557 576
rect 2578 566 2581 643
rect 2578 563 2589 566
rect 2562 483 2565 536
rect 2570 523 2573 546
rect 2498 453 2517 456
rect 2530 453 2541 456
rect 2578 453 2581 526
rect 2490 413 2501 416
rect 2506 413 2509 446
rect 2514 403 2517 453
rect 2466 373 2493 376
rect 2490 346 2493 373
rect 2458 316 2461 346
rect 2490 343 2517 346
rect 2490 333 2493 343
rect 2474 323 2485 326
rect 2490 323 2501 326
rect 2474 316 2477 323
rect 2458 313 2477 316
rect 2506 313 2509 336
rect 2450 303 2461 306
rect 2458 236 2461 303
rect 2458 233 2469 236
rect 2442 213 2453 216
rect 2442 133 2445 213
rect 2458 183 2461 216
rect 2466 133 2469 233
rect 2474 213 2477 276
rect 2514 203 2517 343
rect 2522 213 2525 426
rect 2530 413 2533 436
rect 2538 403 2541 453
rect 2562 413 2565 426
rect 2586 406 2589 563
rect 2562 403 2589 406
rect 2538 226 2541 346
rect 2554 323 2557 346
rect 2562 333 2565 403
rect 2594 386 2597 636
rect 2602 623 2605 693
rect 2634 653 2637 736
rect 2642 646 2645 846
rect 2650 733 2653 903
rect 2658 766 2661 896
rect 2670 836 2673 903
rect 2666 833 2673 836
rect 2666 783 2669 833
rect 2674 803 2677 816
rect 2658 763 2665 766
rect 2650 683 2653 726
rect 2662 676 2665 763
rect 2682 746 2685 933
rect 2634 643 2645 646
rect 2658 673 2665 676
rect 2674 743 2685 746
rect 2610 516 2613 616
rect 2626 543 2629 626
rect 2634 603 2637 643
rect 2606 513 2613 516
rect 2606 436 2609 513
rect 2626 506 2629 536
rect 2634 533 2637 566
rect 2622 503 2629 506
rect 2622 446 2625 503
rect 2538 223 2545 226
rect 2530 183 2533 206
rect 2542 166 2545 223
rect 2554 213 2557 266
rect 2562 223 2565 326
rect 2570 296 2573 386
rect 2590 383 2597 386
rect 2602 433 2609 436
rect 2618 443 2625 446
rect 2578 313 2581 366
rect 2590 296 2593 383
rect 2602 303 2605 433
rect 2618 416 2621 443
rect 2610 413 2621 416
rect 2626 413 2629 436
rect 2610 383 2613 406
rect 2634 403 2637 526
rect 2642 513 2645 606
rect 2650 533 2653 566
rect 2658 486 2661 673
rect 2674 646 2677 743
rect 2682 716 2685 736
rect 2690 733 2693 1116
rect 2698 1033 2701 1126
rect 2706 1026 2709 1153
rect 2698 1023 2709 1026
rect 2698 803 2701 1023
rect 2706 903 2709 966
rect 2714 883 2717 1206
rect 2722 1163 2725 1376
rect 2738 1356 2741 1406
rect 2746 1403 2749 1506
rect 2730 1353 2741 1356
rect 2730 1333 2733 1353
rect 2754 1346 2757 1623
rect 2770 1613 2773 1793
rect 2778 1606 2781 1736
rect 2786 1706 2789 1736
rect 2794 1733 2797 1833
rect 2802 1823 2805 1843
rect 2810 1823 2813 2006
rect 2818 2003 2821 2093
rect 2826 2013 2829 2076
rect 2818 1933 2821 1976
rect 2834 1956 2837 2143
rect 2842 2106 2845 2126
rect 2842 2103 2849 2106
rect 2846 2046 2849 2103
rect 2858 2053 2861 2136
rect 2874 2093 2877 2143
rect 2882 2133 2885 2146
rect 2890 2066 2893 2156
rect 2882 2063 2893 2066
rect 2842 2043 2849 2046
rect 2842 2026 2845 2043
rect 2842 2023 2869 2026
rect 2842 1983 2845 2023
rect 2826 1953 2837 1956
rect 2826 1933 2829 1953
rect 2834 1936 2837 1946
rect 2834 1933 2845 1936
rect 2802 1743 2805 1816
rect 2810 1763 2813 1816
rect 2818 1803 2821 1886
rect 2794 1723 2805 1726
rect 2810 1723 2813 1756
rect 2786 1703 2793 1706
rect 2790 1646 2793 1703
rect 2802 1686 2805 1723
rect 2818 1713 2821 1736
rect 2826 1733 2829 1926
rect 2834 1883 2837 1926
rect 2826 1706 2829 1726
rect 2834 1713 2837 1876
rect 2842 1813 2845 1926
rect 2850 1923 2853 2016
rect 2866 2013 2869 2023
rect 2858 1983 2861 2006
rect 2866 2003 2877 2006
rect 2850 1873 2853 1916
rect 2858 1893 2861 1936
rect 2866 1903 2869 2003
rect 2882 1933 2885 2063
rect 2890 2013 2893 2056
rect 2874 1923 2885 1926
rect 2874 1863 2877 1923
rect 2850 1816 2853 1846
rect 2858 1823 2877 1826
rect 2850 1813 2861 1816
rect 2850 1756 2853 1813
rect 2842 1753 2853 1756
rect 2842 1733 2845 1753
rect 2858 1746 2861 1806
rect 2850 1743 2861 1746
rect 2826 1703 2837 1706
rect 2802 1683 2821 1686
rect 2766 1603 2781 1606
rect 2786 1643 2793 1646
rect 2786 1603 2789 1643
rect 2818 1633 2821 1666
rect 2794 1623 2821 1626
rect 2794 1613 2797 1623
rect 2794 1603 2805 1606
rect 2766 1356 2769 1603
rect 2778 1406 2781 1556
rect 2786 1486 2789 1576
rect 2794 1493 2797 1603
rect 2802 1543 2805 1596
rect 2810 1536 2813 1616
rect 2802 1533 2813 1536
rect 2818 1533 2821 1623
rect 2802 1523 2821 1526
rect 2786 1483 2793 1486
rect 2790 1426 2793 1483
rect 2790 1423 2797 1426
rect 2778 1403 2789 1406
rect 2778 1373 2781 1396
rect 2738 1343 2757 1346
rect 2762 1353 2769 1356
rect 2730 1313 2733 1326
rect 2722 1103 2725 1116
rect 2722 933 2725 1026
rect 2730 1003 2733 1246
rect 2722 873 2725 926
rect 2714 806 2717 816
rect 2706 803 2717 806
rect 2722 803 2725 816
rect 2682 713 2693 716
rect 2706 713 2709 803
rect 2722 776 2725 796
rect 2718 773 2725 776
rect 2670 643 2677 646
rect 2670 596 2673 643
rect 2690 636 2693 713
rect 2718 706 2721 773
rect 2718 703 2725 706
rect 2682 633 2693 636
rect 2682 603 2685 633
rect 2690 596 2693 616
rect 2706 613 2709 636
rect 2670 593 2677 596
rect 2690 593 2697 596
rect 2714 593 2717 686
rect 2674 573 2677 593
rect 2666 513 2669 546
rect 2682 523 2685 556
rect 2694 536 2697 593
rect 2706 536 2709 556
rect 2694 533 2701 536
rect 2706 533 2713 536
rect 2722 533 2725 703
rect 2690 513 2693 526
rect 2658 483 2669 486
rect 2642 413 2645 476
rect 2666 396 2669 483
rect 2698 456 2701 533
rect 2682 453 2701 456
rect 2682 403 2685 453
rect 2710 436 2713 533
rect 2730 526 2733 986
rect 2738 916 2741 1343
rect 2762 1326 2765 1353
rect 2746 1223 2749 1326
rect 2758 1323 2765 1326
rect 2770 1323 2773 1336
rect 2758 1236 2761 1323
rect 2770 1303 2773 1316
rect 2778 1263 2781 1336
rect 2758 1233 2765 1236
rect 2746 1123 2749 1196
rect 2754 1163 2757 1216
rect 2746 963 2749 1086
rect 2754 1013 2757 1066
rect 2762 1033 2765 1233
rect 2770 1223 2773 1256
rect 2770 1173 2773 1216
rect 2778 1203 2781 1226
rect 2786 1193 2789 1403
rect 2762 993 2765 1026
rect 2770 993 2773 1166
rect 2794 1153 2797 1423
rect 2786 1136 2789 1146
rect 2802 1143 2805 1523
rect 2810 1403 2813 1426
rect 2818 1386 2821 1516
rect 2826 1396 2829 1696
rect 2834 1453 2837 1703
rect 2842 1533 2845 1726
rect 2850 1723 2853 1743
rect 2850 1623 2853 1686
rect 2858 1656 2861 1736
rect 2866 1723 2869 1806
rect 2874 1743 2877 1823
rect 2858 1653 2869 1656
rect 2858 1573 2861 1646
rect 2866 1583 2869 1653
rect 2874 1546 2877 1736
rect 2882 1723 2885 1916
rect 2890 1903 2893 1966
rect 2882 1643 2885 1716
rect 2890 1626 2893 1846
rect 2850 1543 2877 1546
rect 2882 1623 2893 1626
rect 2882 1543 2885 1623
rect 2850 1516 2853 1543
rect 2846 1513 2853 1516
rect 2846 1436 2849 1513
rect 2846 1433 2853 1436
rect 2834 1403 2837 1416
rect 2826 1393 2837 1396
rect 2818 1383 2829 1386
rect 2810 1313 2813 1326
rect 2826 1313 2829 1383
rect 2818 1216 2821 1226
rect 2810 1203 2813 1216
rect 2818 1213 2829 1216
rect 2778 1113 2781 1136
rect 2786 1133 2805 1136
rect 2778 1083 2781 1106
rect 2778 983 2781 1006
rect 2786 976 2789 1126
rect 2794 1113 2805 1116
rect 2794 1073 2797 1113
rect 2778 973 2789 976
rect 2746 943 2773 946
rect 2746 923 2749 936
rect 2738 913 2749 916
rect 2738 786 2741 906
rect 2746 806 2749 913
rect 2754 883 2757 936
rect 2746 803 2757 806
rect 2762 803 2765 936
rect 2770 903 2773 943
rect 2778 933 2781 973
rect 2770 803 2773 896
rect 2738 783 2745 786
rect 2742 706 2745 783
rect 2738 703 2745 706
rect 2738 683 2741 703
rect 2754 666 2757 803
rect 2778 796 2781 926
rect 2738 663 2757 666
rect 2762 793 2781 796
rect 2786 796 2789 966
rect 2794 906 2797 1036
rect 2802 943 2805 1106
rect 2810 1023 2813 1156
rect 2818 1093 2821 1126
rect 2826 1003 2829 1196
rect 2834 1013 2837 1393
rect 2842 1253 2845 1416
rect 2850 1383 2853 1433
rect 2850 1323 2853 1336
rect 2858 1306 2861 1536
rect 2890 1533 2893 1616
rect 2898 1613 2901 2376
rect 2906 2236 2909 2436
rect 2914 2256 2917 2426
rect 2922 2393 2925 2416
rect 2938 2413 2941 2426
rect 2946 2416 2949 2513
rect 2978 2506 2981 2553
rect 3026 2546 3029 2613
rect 3034 2586 3037 2606
rect 3042 2593 3053 2596
rect 3034 2583 3045 2586
rect 3026 2543 3033 2546
rect 2978 2503 2989 2506
rect 2954 2423 2981 2426
rect 2946 2413 2957 2416
rect 2930 2353 2933 2406
rect 2954 2403 2957 2413
rect 2938 2333 2949 2336
rect 2954 2326 2957 2396
rect 2962 2386 2965 2416
rect 2978 2403 2981 2423
rect 2986 2403 2989 2503
rect 3002 2426 3005 2536
rect 2998 2423 3005 2426
rect 2962 2383 2981 2386
rect 2922 2303 2925 2326
rect 2930 2323 2957 2326
rect 2962 2316 2965 2356
rect 2970 2333 2973 2366
rect 2978 2323 2981 2383
rect 2986 2373 2989 2396
rect 2998 2366 3001 2423
rect 3010 2393 3013 2416
rect 3018 2373 3021 2496
rect 3030 2426 3033 2543
rect 3030 2423 3037 2426
rect 2998 2363 3005 2366
rect 2962 2313 2969 2316
rect 2914 2253 2941 2256
rect 2906 2233 2917 2236
rect 2906 2193 2909 2216
rect 2914 2213 2917 2233
rect 2914 2133 2917 2146
rect 2906 2013 2909 2126
rect 2922 2046 2925 2166
rect 2930 2113 2933 2126
rect 2938 2103 2941 2253
rect 2918 2043 2925 2046
rect 2906 1823 2909 2006
rect 2918 1956 2921 2043
rect 2930 2003 2933 2036
rect 2938 2013 2941 2026
rect 2938 1983 2941 1996
rect 2918 1953 2925 1956
rect 2914 1833 2917 1936
rect 2914 1806 2917 1826
rect 2906 1803 2917 1806
rect 2906 1556 2909 1746
rect 2914 1733 2917 1776
rect 2914 1623 2917 1646
rect 2914 1603 2917 1616
rect 2898 1553 2909 1556
rect 2866 1523 2885 1526
rect 2898 1523 2901 1553
rect 2866 1406 2869 1446
rect 2866 1403 2877 1406
rect 2866 1333 2869 1396
rect 2874 1386 2877 1403
rect 2882 1393 2885 1446
rect 2874 1383 2885 1386
rect 2854 1303 2861 1306
rect 2842 1093 2845 1246
rect 2854 1236 2857 1303
rect 2854 1233 2861 1236
rect 2850 1173 2853 1216
rect 2850 1123 2853 1136
rect 2858 1106 2861 1233
rect 2866 1203 2869 1316
rect 2866 1143 2869 1196
rect 2854 1103 2861 1106
rect 2854 1026 2857 1103
rect 2802 923 2805 936
rect 2794 903 2801 906
rect 2798 806 2801 903
rect 2810 823 2813 986
rect 2818 923 2821 956
rect 2834 913 2837 946
rect 2818 826 2821 876
rect 2826 833 2829 906
rect 2818 823 2829 826
rect 2810 813 2821 816
rect 2798 803 2821 806
rect 2786 793 2797 796
rect 2738 603 2741 663
rect 2754 613 2757 656
rect 2746 553 2749 606
rect 2746 526 2749 536
rect 2754 533 2757 606
rect 2762 586 2765 793
rect 2770 603 2773 726
rect 2762 583 2769 586
rect 2698 423 2701 436
rect 2706 433 2713 436
rect 2722 523 2733 526
rect 2738 523 2749 526
rect 2706 416 2709 433
rect 2698 413 2709 416
rect 2722 416 2725 523
rect 2730 423 2733 466
rect 2722 413 2733 416
rect 2666 393 2673 396
rect 2626 333 2645 336
rect 2650 333 2653 346
rect 2658 333 2661 386
rect 2642 326 2645 333
rect 2634 306 2637 326
rect 2642 323 2653 326
rect 2670 316 2673 393
rect 2682 323 2685 336
rect 2698 333 2701 413
rect 2626 303 2637 306
rect 2570 293 2581 296
rect 2590 293 2597 296
rect 2554 173 2557 206
rect 2542 163 2549 166
rect 2410 63 2413 126
rect 2498 103 2501 156
rect 2530 123 2533 136
rect 2546 113 2549 163
rect 2554 93 2557 106
rect 2562 63 2565 206
rect 2578 136 2581 293
rect 2594 276 2597 293
rect 2594 273 2605 276
rect 2602 226 2605 273
rect 2626 236 2629 303
rect 2650 243 2653 316
rect 2666 313 2673 316
rect 2706 313 2709 406
rect 2738 396 2741 523
rect 2746 443 2749 516
rect 2754 513 2757 526
rect 2766 516 2769 583
rect 2778 533 2781 746
rect 2794 706 2797 793
rect 2786 703 2797 706
rect 2786 603 2789 703
rect 2794 603 2797 696
rect 2802 606 2805 736
rect 2810 683 2813 746
rect 2810 613 2813 646
rect 2802 603 2813 606
rect 2810 593 2813 603
rect 2818 576 2821 803
rect 2826 726 2829 823
rect 2834 763 2837 826
rect 2842 733 2845 1026
rect 2854 1023 2861 1026
rect 2850 993 2853 1006
rect 2850 733 2853 926
rect 2858 893 2861 1023
rect 2866 913 2869 1136
rect 2874 1106 2877 1376
rect 2882 1303 2885 1383
rect 2890 1343 2893 1516
rect 2906 1433 2909 1546
rect 2914 1523 2917 1536
rect 2922 1473 2925 1953
rect 2930 1923 2933 1966
rect 2938 1943 2941 1956
rect 2938 1923 2941 1936
rect 2930 1603 2933 1916
rect 2938 1783 2941 1826
rect 2938 1733 2941 1756
rect 2946 1656 2949 2266
rect 2954 2213 2957 2296
rect 2966 2246 2969 2313
rect 3002 2256 3005 2363
rect 3026 2323 3029 2416
rect 3034 2316 3037 2423
rect 2962 2243 2969 2246
rect 2978 2253 3005 2256
rect 3026 2313 3037 2316
rect 3042 2313 3045 2583
rect 3074 2543 3077 2606
rect 3086 2546 3089 2623
rect 3106 2616 3109 2653
rect 3098 2613 3109 2616
rect 3114 2613 3117 2646
rect 3086 2543 3093 2546
rect 3050 2523 3053 2536
rect 3082 2506 3085 2526
rect 3074 2503 3085 2506
rect 3074 2446 3077 2503
rect 3090 2493 3093 2543
rect 3066 2443 3077 2446
rect 3050 2413 3053 2426
rect 3050 2323 3053 2396
rect 2954 2013 2957 2116
rect 2962 2096 2965 2243
rect 2978 2203 2981 2253
rect 3026 2243 3029 2313
rect 3026 2213 3029 2226
rect 2978 2133 2981 2196
rect 3058 2143 3061 2216
rect 3066 2213 3069 2443
rect 3090 2436 3093 2486
rect 3082 2433 3093 2436
rect 3082 2406 3085 2433
rect 3090 2413 3093 2426
rect 3074 2403 3085 2406
rect 3098 2403 3101 2566
rect 3106 2553 3109 2606
rect 3114 2523 3117 2606
rect 3122 2526 3125 2653
rect 3134 2586 3137 2663
rect 3130 2583 3137 2586
rect 3146 2623 3181 2626
rect 3130 2533 3133 2583
rect 3138 2533 3141 2566
rect 3122 2523 3141 2526
rect 3146 2523 3149 2623
rect 3154 2543 3157 2606
rect 3162 2546 3165 2616
rect 3178 2613 3181 2623
rect 3170 2553 3173 2606
rect 3178 2593 3181 2606
rect 3162 2543 3173 2546
rect 3154 2533 3165 2536
rect 3154 2523 3165 2526
rect 3106 2513 3133 2516
rect 3106 2496 3109 2513
rect 3138 2506 3141 2523
rect 3170 2513 3173 2543
rect 3178 2523 3181 2536
rect 3186 2506 3189 2726
rect 3198 2636 3201 2733
rect 3230 2716 3233 2763
rect 3250 2743 3253 2803
rect 3290 2793 3293 2803
rect 3298 2766 3301 2806
rect 3306 2793 3309 2813
rect 3290 2763 3301 2766
rect 3242 2733 3253 2736
rect 3242 2723 3245 2733
rect 3230 2713 3237 2716
rect 3130 2503 3141 2506
rect 3182 2503 3189 2506
rect 3194 2633 3201 2636
rect 3106 2493 3117 2496
rect 3114 2436 3117 2493
rect 3106 2433 3117 2436
rect 3106 2413 3109 2433
rect 3130 2423 3133 2503
rect 3182 2436 3185 2503
rect 3182 2433 3189 2436
rect 3138 2423 3173 2426
rect 3114 2413 3133 2416
rect 3026 2113 3029 2126
rect 2962 2093 2969 2096
rect 2966 2026 2969 2093
rect 2962 2023 2969 2026
rect 2954 1933 2957 1976
rect 2954 1903 2957 1926
rect 2954 1813 2957 1836
rect 2954 1753 2957 1806
rect 2954 1733 2957 1746
rect 2954 1713 2957 1726
rect 2938 1653 2949 1656
rect 2938 1613 2941 1653
rect 2930 1523 2933 1576
rect 2938 1533 2941 1566
rect 2898 1403 2901 1426
rect 2890 1286 2893 1316
rect 2886 1283 2893 1286
rect 2886 1216 2889 1283
rect 2882 1213 2889 1216
rect 2882 1193 2885 1213
rect 2898 1206 2901 1396
rect 2906 1393 2909 1406
rect 2914 1346 2917 1466
rect 2906 1343 2917 1346
rect 2906 1243 2909 1343
rect 2914 1323 2917 1336
rect 2922 1236 2925 1436
rect 2930 1416 2933 1456
rect 2938 1423 2941 1516
rect 2930 1413 2941 1416
rect 2930 1326 2933 1396
rect 2938 1373 2941 1413
rect 2938 1333 2941 1346
rect 2930 1323 2941 1326
rect 2938 1303 2941 1316
rect 2890 1203 2901 1206
rect 2906 1233 2925 1236
rect 2890 1186 2893 1203
rect 2882 1183 2893 1186
rect 2882 1123 2885 1183
rect 2874 1103 2881 1106
rect 2890 1103 2893 1146
rect 2898 1123 2901 1196
rect 2906 1143 2909 1233
rect 2922 1223 2933 1226
rect 2878 1026 2881 1103
rect 2878 1023 2885 1026
rect 2874 906 2877 1016
rect 2882 923 2885 1023
rect 2866 903 2877 906
rect 2882 903 2885 916
rect 2826 723 2853 726
rect 2826 703 2829 716
rect 2858 713 2861 826
rect 2866 813 2869 903
rect 2890 893 2893 1046
rect 2906 1023 2909 1136
rect 2914 1133 2917 1216
rect 2938 1213 2941 1256
rect 2922 1133 2933 1136
rect 2826 603 2829 616
rect 2762 513 2769 516
rect 2762 496 2765 513
rect 2758 493 2765 496
rect 2730 393 2741 396
rect 2666 293 2669 313
rect 2626 233 2637 236
rect 2594 223 2605 226
rect 2594 203 2597 223
rect 2634 213 2637 233
rect 2658 206 2661 216
rect 2634 203 2661 206
rect 2570 133 2581 136
rect 2666 133 2669 226
rect 2570 113 2573 133
rect 2602 63 2605 126
rect 2674 123 2677 206
rect 2682 73 2685 226
rect 2690 103 2693 216
rect 2714 206 2717 326
rect 2730 223 2733 393
rect 2758 386 2761 493
rect 2770 403 2773 486
rect 2786 416 2789 576
rect 2810 573 2821 576
rect 2810 516 2813 573
rect 2834 523 2837 686
rect 2842 603 2845 626
rect 2858 593 2861 656
rect 2874 613 2877 836
rect 2882 823 2885 876
rect 2890 736 2893 826
rect 2882 733 2893 736
rect 2882 723 2885 733
rect 2890 703 2893 716
rect 2858 533 2861 566
rect 2810 513 2853 516
rect 2834 496 2837 513
rect 2782 413 2789 416
rect 2802 426 2805 496
rect 2830 493 2837 496
rect 2802 423 2821 426
rect 2758 383 2765 386
rect 2762 363 2765 383
rect 2782 356 2785 413
rect 2794 393 2797 406
rect 2802 403 2805 423
rect 2810 363 2813 416
rect 2818 413 2821 423
rect 2830 396 2833 493
rect 2858 466 2861 526
rect 2866 493 2869 606
rect 2890 586 2893 606
rect 2886 583 2893 586
rect 2874 523 2877 576
rect 2886 496 2889 583
rect 2898 516 2901 1016
rect 2914 1003 2917 1126
rect 2922 986 2925 1016
rect 2918 983 2925 986
rect 2918 916 2921 983
rect 2906 723 2909 916
rect 2914 913 2921 916
rect 2930 913 2933 1056
rect 2906 653 2909 716
rect 2906 536 2909 646
rect 2914 603 2917 913
rect 2922 863 2925 906
rect 2922 813 2925 826
rect 2922 686 2925 776
rect 2930 733 2933 856
rect 2938 706 2941 1146
rect 2946 1136 2949 1646
rect 2954 1543 2957 1626
rect 2954 1493 2957 1536
rect 2954 1333 2957 1486
rect 2962 1396 2965 2023
rect 2970 1983 2973 2006
rect 2970 1923 2973 1956
rect 2970 1773 2973 1896
rect 2970 1723 2973 1756
rect 2970 1533 2973 1616
rect 2970 1513 2973 1526
rect 2970 1413 2973 1476
rect 2978 1466 2981 2066
rect 2986 1913 2989 2036
rect 2994 1826 2997 2026
rect 3002 2013 3013 2016
rect 3026 2006 3029 2046
rect 3002 2003 3029 2006
rect 3002 1843 3005 2003
rect 3042 1986 3045 2136
rect 3066 2123 3069 2206
rect 3074 2133 3077 2403
rect 3114 2386 3117 2413
rect 3122 2403 3133 2406
rect 3122 2393 3125 2403
rect 3138 2396 3141 2423
rect 3154 2406 3157 2416
rect 3186 2413 3189 2433
rect 3130 2393 3141 2396
rect 3082 2106 3085 2386
rect 3114 2383 3125 2386
rect 3074 2103 3085 2106
rect 3074 2056 3077 2103
rect 3074 2053 3085 2056
rect 3082 2033 3085 2053
rect 3058 2023 3085 2026
rect 3058 2013 3061 2023
rect 3050 1993 3053 2006
rect 3066 1986 3069 2016
rect 3034 1983 3069 1986
rect 2994 1823 3005 1826
rect 2986 1813 2997 1816
rect 2986 1763 2989 1806
rect 2994 1783 2997 1806
rect 2994 1746 2997 1776
rect 2990 1743 2997 1746
rect 2990 1626 2993 1743
rect 2990 1623 2997 1626
rect 2986 1563 2989 1606
rect 2994 1603 2997 1623
rect 3002 1573 3005 1823
rect 3010 1733 3013 1976
rect 3018 1873 3021 1936
rect 3026 1923 3029 1956
rect 3034 1883 3037 1983
rect 3018 1723 3021 1806
rect 3026 1763 3029 1826
rect 3026 1703 3029 1736
rect 3034 1723 3037 1806
rect 3042 1673 3045 1936
rect 3050 1763 3053 1926
rect 3058 1923 3069 1926
rect 3050 1733 3053 1746
rect 3010 1603 3013 1666
rect 2986 1533 2997 1536
rect 3002 1526 3005 1536
rect 2986 1483 2989 1526
rect 2994 1523 3005 1526
rect 3010 1523 3013 1536
rect 2978 1463 2985 1466
rect 2982 1406 2985 1463
rect 2978 1403 2985 1406
rect 2962 1393 2969 1396
rect 2954 1213 2957 1316
rect 2966 1246 2969 1393
rect 2962 1243 2969 1246
rect 2954 1153 2957 1206
rect 2946 1133 2953 1136
rect 2950 1066 2953 1133
rect 2946 1063 2953 1066
rect 2946 1043 2949 1063
rect 2946 1013 2949 1036
rect 2954 1003 2957 1026
rect 2962 1013 2965 1243
rect 2970 1203 2973 1226
rect 2970 1013 2973 1136
rect 2946 823 2949 956
rect 2954 936 2957 946
rect 2954 933 2965 936
rect 2954 823 2957 926
rect 2962 816 2965 933
rect 2946 803 2949 816
rect 2954 813 2965 816
rect 2954 716 2957 813
rect 2946 713 2957 716
rect 2938 703 2949 706
rect 2922 683 2933 686
rect 2930 626 2933 683
rect 2922 623 2933 626
rect 2922 596 2925 623
rect 2914 593 2925 596
rect 2914 546 2917 593
rect 2938 563 2941 606
rect 2914 543 2933 546
rect 2906 533 2925 536
rect 2922 516 2925 533
rect 2930 526 2933 543
rect 2938 533 2941 546
rect 2930 523 2941 526
rect 2946 523 2949 703
rect 2954 613 2957 626
rect 2954 583 2957 606
rect 2954 533 2957 576
rect 2962 536 2965 746
rect 2970 556 2973 1006
rect 2978 943 2981 1403
rect 2994 1386 2997 1523
rect 3018 1516 3021 1616
rect 3026 1613 3045 1616
rect 3026 1593 3029 1606
rect 3034 1553 3037 1576
rect 3034 1533 3037 1546
rect 3042 1533 3045 1606
rect 3010 1513 3021 1516
rect 2990 1383 2997 1386
rect 2990 1326 2993 1383
rect 3002 1343 3005 1486
rect 3010 1393 3013 1513
rect 2990 1323 2997 1326
rect 2986 1186 2989 1306
rect 2994 1253 2997 1323
rect 2994 1196 2997 1216
rect 3002 1206 3005 1336
rect 3018 1326 3021 1506
rect 3026 1333 3029 1516
rect 3034 1413 3037 1516
rect 3042 1423 3045 1436
rect 3010 1306 3013 1326
rect 3018 1323 3029 1326
rect 3010 1303 3017 1306
rect 3014 1236 3017 1303
rect 3014 1233 3021 1236
rect 3002 1203 3013 1206
rect 2994 1193 3005 1196
rect 2986 1183 2997 1186
rect 2986 933 2989 1176
rect 2994 1106 2997 1183
rect 3002 1123 3005 1193
rect 2994 1103 3001 1106
rect 2998 1026 3001 1103
rect 3010 1033 3013 1116
rect 3018 1103 3021 1233
rect 3026 1223 3029 1323
rect 3026 1036 3029 1216
rect 3034 1203 3037 1326
rect 3042 1303 3045 1356
rect 3042 1203 3045 1286
rect 3034 1123 3037 1146
rect 3026 1033 3033 1036
rect 2998 1023 3021 1026
rect 2994 986 2997 1016
rect 3002 1003 3005 1016
rect 2994 983 3001 986
rect 2998 926 3001 983
rect 2994 923 3001 926
rect 2978 803 2981 866
rect 2978 703 2981 796
rect 2986 723 2989 816
rect 2978 563 2981 616
rect 2994 603 2997 923
rect 3002 833 3005 866
rect 3002 793 3005 826
rect 3010 823 3013 926
rect 3018 913 3021 1023
rect 3030 956 3033 1033
rect 3026 953 3033 956
rect 3018 816 3021 836
rect 3010 813 3021 816
rect 3002 713 3005 726
rect 3010 696 3013 806
rect 3006 693 3013 696
rect 3006 556 3009 693
rect 3018 566 3021 786
rect 3026 773 3029 953
rect 3026 633 3029 766
rect 3018 563 3025 566
rect 2970 553 2981 556
rect 3006 553 3013 556
rect 2962 533 2973 536
rect 2978 533 2981 553
rect 2898 513 2909 516
rect 2886 493 2893 496
rect 2826 393 2833 396
rect 2842 463 2861 466
rect 2782 353 2789 356
rect 2738 333 2781 336
rect 2762 323 2773 326
rect 2754 303 2757 316
rect 2706 203 2717 206
rect 2730 123 2733 206
rect 2746 203 2749 216
rect 2762 213 2765 316
rect 2778 313 2781 333
rect 2786 306 2789 353
rect 2826 346 2829 393
rect 2770 303 2789 306
rect 2738 123 2741 136
rect 2746 133 2757 136
rect 2314 33 2317 63
rect 2770 13 2773 296
rect 2786 133 2789 276
rect 2794 196 2797 346
rect 2826 343 2837 346
rect 2802 313 2805 336
rect 2834 326 2837 343
rect 2842 336 2845 463
rect 2850 396 2853 416
rect 2850 393 2885 396
rect 2842 333 2853 336
rect 2834 323 2845 326
rect 2850 306 2853 333
rect 2858 313 2861 386
rect 2866 323 2869 336
rect 2842 303 2853 306
rect 2874 303 2877 326
rect 2842 246 2845 303
rect 2842 243 2853 246
rect 2802 223 2845 226
rect 2802 203 2805 223
rect 2818 203 2821 216
rect 2794 193 2813 196
rect 2794 113 2797 166
rect 2810 136 2813 193
rect 2810 133 2821 136
rect 2818 63 2821 126
rect 2826 113 2829 216
rect 2842 213 2845 223
rect 2834 183 2837 206
rect 2850 203 2853 243
rect 2866 193 2869 296
rect 2882 253 2885 393
rect 2890 343 2893 493
rect 2906 436 2909 513
rect 2898 433 2909 436
rect 2918 513 2925 516
rect 2882 176 2885 206
rect 2890 183 2893 326
rect 2898 273 2901 433
rect 2918 426 2921 513
rect 2918 423 2925 426
rect 2906 403 2909 416
rect 2906 263 2909 396
rect 2914 203 2917 406
rect 2922 176 2925 423
rect 2858 113 2861 126
rect 2866 113 2869 136
rect 2874 123 2877 176
rect 2882 173 2925 176
rect 2882 156 2885 173
rect 2930 156 2933 516
rect 2938 506 2941 523
rect 2938 503 2957 506
rect 2946 413 2949 436
rect 2954 413 2957 503
rect 2962 496 2965 526
rect 2970 513 2973 533
rect 2986 523 2989 546
rect 3002 506 3005 536
rect 2994 503 3005 506
rect 2962 493 2973 496
rect 2970 426 2973 493
rect 2994 456 2997 503
rect 2994 453 3005 456
rect 2962 423 2973 426
rect 2962 396 2965 423
rect 2954 393 2965 396
rect 2954 336 2957 393
rect 2970 353 2973 406
rect 2954 333 2965 336
rect 2938 296 2941 326
rect 2938 293 2949 296
rect 2946 246 2949 293
rect 2962 283 2965 333
rect 2970 293 2973 326
rect 2994 306 2997 416
rect 3002 403 3005 453
rect 2978 303 2997 306
rect 2942 243 2949 246
rect 2942 166 2945 243
rect 2954 223 2989 226
rect 2954 213 2957 223
rect 2962 203 2965 216
rect 2970 176 2973 206
rect 2978 203 2981 216
rect 2986 203 2989 223
rect 2970 173 2989 176
rect 2994 173 2997 216
rect 2882 153 2893 156
rect 2890 106 2893 153
rect 2882 103 2893 106
rect 2922 153 2933 156
rect 2938 163 2945 166
rect 2882 33 2885 103
rect 2922 76 2925 153
rect 2938 83 2941 163
rect 2946 133 2949 146
rect 2970 133 2973 166
rect 2986 136 2989 173
rect 2978 126 2981 136
rect 2986 133 2997 136
rect 3002 126 3005 316
rect 2954 123 2973 126
rect 2978 123 3005 126
rect 2970 103 2973 116
rect 3010 113 3013 553
rect 3022 486 3025 563
rect 3018 483 3025 486
rect 3018 463 3021 483
rect 3018 423 3021 436
rect 3034 406 3037 936
rect 3042 873 3045 1186
rect 3050 1013 3053 1716
rect 3058 1713 3061 1856
rect 3066 1803 3069 1923
rect 3074 1793 3077 1986
rect 3082 1933 3085 2006
rect 3082 1823 3085 1856
rect 3082 1783 3085 1806
rect 3074 1733 3077 1776
rect 3058 1603 3061 1706
rect 3066 1623 3069 1686
rect 3058 1353 3061 1536
rect 3066 1513 3069 1616
rect 3074 1543 3077 1726
rect 3082 1623 3085 1766
rect 3090 1716 3093 2306
rect 3114 2273 3117 2336
rect 3122 2296 3125 2383
rect 3130 2323 3133 2393
rect 3146 2343 3149 2406
rect 3154 2403 3189 2406
rect 3138 2333 3157 2336
rect 3130 2303 3133 2316
rect 3138 2296 3141 2326
rect 3122 2293 3141 2296
rect 3098 2213 3101 2246
rect 3122 2213 3125 2226
rect 3130 2166 3133 2216
rect 3122 2163 3133 2166
rect 3122 2156 3125 2163
rect 3098 2153 3125 2156
rect 3098 2123 3101 2153
rect 3106 2113 3109 2136
rect 3122 2133 3125 2146
rect 3130 2133 3133 2156
rect 3114 2123 3125 2126
rect 3138 2123 3141 2196
rect 3154 2146 3157 2333
rect 3170 2316 3173 2396
rect 3186 2333 3189 2396
rect 3166 2313 3173 2316
rect 3166 2246 3169 2313
rect 3166 2243 3173 2246
rect 3162 2213 3165 2226
rect 3154 2143 3165 2146
rect 3146 2133 3157 2136
rect 3098 2003 3101 2026
rect 3106 1976 3109 2016
rect 3098 1973 3109 1976
rect 3098 1913 3101 1973
rect 3106 1933 3109 1966
rect 3114 1916 3117 2106
rect 3122 2093 3125 2123
rect 3154 2093 3157 2126
rect 3162 2053 3165 2143
rect 3154 2006 3157 2016
rect 3110 1913 3117 1916
rect 3122 2003 3157 2006
rect 3110 1846 3113 1913
rect 3110 1843 3117 1846
rect 3106 1816 3109 1826
rect 3098 1813 3109 1816
rect 3098 1753 3101 1813
rect 3106 1773 3109 1806
rect 3090 1713 3101 1716
rect 3090 1643 3093 1713
rect 3098 1626 3101 1706
rect 3090 1623 3101 1626
rect 3066 1403 3069 1416
rect 3074 1403 3077 1536
rect 3082 1413 3085 1616
rect 3090 1613 3093 1623
rect 3090 1543 3093 1606
rect 3090 1483 3093 1526
rect 3098 1466 3101 1616
rect 3106 1543 3109 1766
rect 3114 1743 3117 1843
rect 3114 1703 3117 1736
rect 3114 1603 3117 1636
rect 3094 1463 3101 1466
rect 3094 1366 3097 1463
rect 3106 1443 3109 1536
rect 3114 1506 3117 1586
rect 3122 1533 3125 2003
rect 3146 1993 3157 1996
rect 3162 1986 3165 2046
rect 3154 1983 3165 1986
rect 3130 1943 3141 1946
rect 3130 1903 3133 1926
rect 3138 1913 3141 1926
rect 3146 1853 3149 1976
rect 3154 1913 3157 1983
rect 3162 1943 3165 1956
rect 3170 1936 3173 2243
rect 3178 2213 3181 2306
rect 3186 2303 3189 2316
rect 3178 2156 3181 2206
rect 3186 2203 3189 2236
rect 3194 2163 3197 2633
rect 3202 2516 3205 2616
rect 3210 2533 3213 2696
rect 3218 2616 3221 2636
rect 3218 2613 3225 2616
rect 3222 2546 3225 2613
rect 3218 2543 3225 2546
rect 3202 2513 3209 2516
rect 3206 2456 3209 2513
rect 3218 2506 3221 2543
rect 3234 2526 3237 2713
rect 3274 2706 3277 2726
rect 3266 2703 3277 2706
rect 3266 2656 3269 2703
rect 3266 2653 3277 2656
rect 3274 2633 3277 2653
rect 3282 2626 3285 2726
rect 3290 2723 3293 2763
rect 3322 2736 3325 2806
rect 3346 2796 3349 2806
rect 3370 2803 3381 2806
rect 3346 2793 3365 2796
rect 3322 2733 3341 2736
rect 3306 2693 3309 2716
rect 3314 2703 3317 2726
rect 3322 2703 3325 2733
rect 3330 2636 3333 2716
rect 3346 2706 3349 2726
rect 3342 2703 3349 2706
rect 3342 2646 3345 2703
rect 3342 2643 3349 2646
rect 3250 2623 3285 2626
rect 3306 2633 3333 2636
rect 3242 2533 3245 2606
rect 3250 2593 3253 2623
rect 3266 2613 3293 2616
rect 3258 2546 3261 2606
rect 3274 2583 3277 2606
rect 3282 2576 3285 2606
rect 3274 2573 3285 2576
rect 3250 2543 3261 2546
rect 3266 2533 3269 2546
rect 3234 2523 3265 2526
rect 3218 2503 3237 2506
rect 3206 2453 3221 2456
rect 3202 2366 3205 2416
rect 3218 2413 3221 2453
rect 3210 2383 3213 2406
rect 3218 2403 3229 2406
rect 3234 2403 3237 2503
rect 3242 2496 3245 2516
rect 3242 2493 3253 2496
rect 3250 2436 3253 2493
rect 3242 2433 3253 2436
rect 3202 2363 3209 2366
rect 3206 2286 3209 2363
rect 3218 2323 3221 2403
rect 3242 2396 3245 2433
rect 3262 2426 3265 2523
rect 3262 2423 3269 2426
rect 3250 2403 3253 2416
rect 3234 2393 3245 2396
rect 3218 2306 3221 2316
rect 3234 2313 3237 2393
rect 3250 2383 3253 2396
rect 3258 2393 3261 2406
rect 3250 2323 3253 2336
rect 3266 2326 3269 2423
rect 3274 2416 3277 2573
rect 3282 2533 3285 2556
rect 3290 2536 3293 2613
rect 3298 2573 3301 2616
rect 3290 2533 3301 2536
rect 3290 2506 3293 2526
rect 3286 2503 3293 2506
rect 3286 2446 3289 2503
rect 3286 2443 3293 2446
rect 3290 2426 3293 2443
rect 3298 2433 3301 2533
rect 3290 2423 3301 2426
rect 3274 2413 3293 2416
rect 3266 2323 3277 2326
rect 3242 2306 3245 2316
rect 3218 2303 3245 2306
rect 3250 2303 3253 2316
rect 3266 2303 3269 2316
rect 3206 2283 3213 2286
rect 3210 2226 3213 2283
rect 3242 2263 3245 2303
rect 3202 2223 3213 2226
rect 3202 2206 3205 2223
rect 3226 2206 3229 2216
rect 3202 2203 3221 2206
rect 3226 2203 3237 2206
rect 3226 2173 3229 2196
rect 3178 2153 3197 2156
rect 3178 1943 3181 2136
rect 3194 2133 3197 2153
rect 3218 2086 3221 2146
rect 3226 2123 3229 2136
rect 3234 2106 3237 2203
rect 3202 2083 3221 2086
rect 3230 2103 3237 2106
rect 3202 2066 3205 2083
rect 3202 2063 3213 2066
rect 3170 1933 3181 1936
rect 3186 1933 3189 2056
rect 3210 2016 3213 2063
rect 3202 2013 3213 2016
rect 3162 1896 3165 1926
rect 3158 1893 3165 1896
rect 3130 1736 3133 1826
rect 3158 1816 3161 1893
rect 3138 1793 3141 1816
rect 3146 1813 3161 1816
rect 3170 1816 3173 1926
rect 3178 1923 3181 1933
rect 3178 1816 3181 1826
rect 3170 1813 3181 1816
rect 3130 1733 3141 1736
rect 3130 1593 3133 1726
rect 3138 1573 3141 1733
rect 3146 1683 3149 1813
rect 3154 1803 3173 1806
rect 3154 1693 3157 1803
rect 3162 1626 3165 1776
rect 3178 1746 3181 1813
rect 3186 1806 3189 1916
rect 3194 1893 3197 1936
rect 3202 1863 3205 2013
rect 3230 2006 3233 2103
rect 3230 2003 3237 2006
rect 3218 1933 3221 1996
rect 3234 1983 3237 2003
rect 3218 1896 3221 1926
rect 3214 1893 3221 1896
rect 3214 1836 3217 1893
rect 3214 1833 3221 1836
rect 3202 1816 3205 1826
rect 3202 1813 3213 1816
rect 3186 1803 3205 1806
rect 3202 1783 3205 1803
rect 3210 1793 3213 1813
rect 3170 1743 3197 1746
rect 3170 1723 3173 1743
rect 3186 1716 3189 1736
rect 3194 1733 3197 1743
rect 3182 1713 3189 1716
rect 3146 1623 3165 1626
rect 3146 1566 3149 1623
rect 3154 1603 3157 1616
rect 3162 1593 3165 1606
rect 3146 1563 3157 1566
rect 3122 1513 3125 1526
rect 3114 1503 3125 1506
rect 3130 1503 3133 1546
rect 3146 1523 3149 1556
rect 3122 1416 3125 1503
rect 3130 1423 3133 1436
rect 3106 1413 3117 1416
rect 3122 1413 3133 1416
rect 3074 1363 3097 1366
rect 3058 1303 3061 1316
rect 3074 1296 3077 1363
rect 3090 1323 3093 1346
rect 3098 1303 3101 1356
rect 3066 1293 3077 1296
rect 3058 1213 3061 1226
rect 3050 923 3053 936
rect 3042 763 3045 836
rect 3050 793 3053 856
rect 3042 706 3045 756
rect 3050 723 3053 786
rect 3042 703 3049 706
rect 3046 626 3049 703
rect 3042 623 3049 626
rect 3042 586 3045 623
rect 3058 613 3061 1206
rect 3066 1043 3069 1293
rect 3106 1286 3109 1406
rect 3114 1323 3117 1413
rect 3102 1283 3109 1286
rect 3066 1023 3069 1036
rect 3066 993 3069 1016
rect 3066 813 3069 976
rect 3074 806 3077 1226
rect 3082 1193 3085 1226
rect 3082 1133 3085 1146
rect 3082 1113 3085 1126
rect 3082 1003 3085 1106
rect 3082 923 3085 996
rect 3066 803 3077 806
rect 3082 803 3085 896
rect 3066 706 3069 803
rect 3090 783 3093 1276
rect 3102 1226 3105 1283
rect 3098 1223 3105 1226
rect 3098 1026 3101 1223
rect 3114 1216 3117 1316
rect 3122 1223 3125 1406
rect 3130 1333 3133 1413
rect 3130 1313 3133 1326
rect 3138 1313 3141 1496
rect 3154 1476 3157 1563
rect 3146 1473 3157 1476
rect 3146 1333 3149 1473
rect 3138 1223 3141 1296
rect 3106 1213 3117 1216
rect 3106 1033 3109 1213
rect 3114 1153 3117 1206
rect 3122 1193 3125 1216
rect 3130 1213 3141 1216
rect 3130 1183 3133 1213
rect 3138 1163 3141 1206
rect 3146 1203 3149 1326
rect 3154 1173 3157 1406
rect 3162 1393 3165 1586
rect 3170 1573 3173 1686
rect 3182 1646 3185 1713
rect 3194 1656 3197 1716
rect 3202 1693 3205 1746
rect 3194 1653 3201 1656
rect 3182 1643 3189 1646
rect 3178 1556 3181 1626
rect 3186 1593 3189 1643
rect 3198 1576 3201 1653
rect 3210 1583 3213 1766
rect 3174 1553 3181 1556
rect 3174 1376 3177 1553
rect 3186 1403 3189 1576
rect 3198 1573 3213 1576
rect 3194 1503 3197 1536
rect 3202 1513 3205 1526
rect 3210 1513 3213 1573
rect 3202 1413 3205 1506
rect 3218 1496 3221 1833
rect 3226 1613 3229 1856
rect 3234 1763 3237 1866
rect 3242 1743 3245 2216
rect 3250 2193 3253 2216
rect 3258 2203 3261 2226
rect 3258 2043 3261 2166
rect 3266 1993 3269 2256
rect 3274 2116 3277 2323
rect 3282 2136 3285 2246
rect 3290 2183 3293 2336
rect 3298 2323 3301 2423
rect 3306 2396 3309 2633
rect 3314 2623 3341 2626
rect 3314 2613 3317 2623
rect 3322 2563 3325 2606
rect 3330 2573 3333 2606
rect 3322 2426 3325 2506
rect 3330 2496 3333 2556
rect 3338 2503 3341 2623
rect 3346 2616 3349 2643
rect 3354 2626 3357 2716
rect 3362 2693 3365 2706
rect 3386 2626 3389 2716
rect 3394 2703 3397 2816
rect 3354 2623 3373 2626
rect 3386 2623 3397 2626
rect 3346 2613 3365 2616
rect 3370 2606 3373 2623
rect 3346 2603 3373 2606
rect 3346 2593 3349 2603
rect 3346 2513 3349 2526
rect 3354 2513 3357 2546
rect 3362 2523 3365 2596
rect 3378 2543 3381 2616
rect 3394 2576 3397 2623
rect 3386 2573 3397 2576
rect 3386 2553 3389 2573
rect 3354 2496 3357 2506
rect 3330 2493 3357 2496
rect 3330 2433 3357 2436
rect 3322 2423 3341 2426
rect 3322 2413 3341 2416
rect 3306 2393 3317 2396
rect 3314 2316 3317 2393
rect 3330 2316 3333 2346
rect 3338 2323 3341 2413
rect 3346 2403 3349 2416
rect 3354 2356 3357 2433
rect 3362 2403 3365 2506
rect 3378 2503 3381 2516
rect 3386 2426 3389 2446
rect 3386 2423 3397 2426
rect 3354 2353 3373 2356
rect 3354 2333 3357 2346
rect 3362 2323 3365 2336
rect 3298 2276 3301 2316
rect 3306 2313 3317 2316
rect 3326 2313 3333 2316
rect 3338 2313 3357 2316
rect 3306 2293 3309 2313
rect 3298 2273 3309 2276
rect 3306 2226 3309 2273
rect 3326 2246 3329 2313
rect 3326 2243 3333 2246
rect 3298 2223 3309 2226
rect 3298 2166 3301 2223
rect 3322 2213 3325 2226
rect 3330 2213 3333 2243
rect 3298 2163 3317 2166
rect 3282 2133 3301 2136
rect 3298 2123 3301 2133
rect 3274 2113 3285 2116
rect 3282 2056 3285 2113
rect 3282 2053 3293 2056
rect 3290 2036 3293 2053
rect 3290 2033 3297 2036
rect 3250 1883 3253 1956
rect 3258 1906 3261 1946
rect 3266 1923 3269 1986
rect 3258 1903 3265 1906
rect 3250 1823 3253 1846
rect 3250 1803 3253 1816
rect 3262 1796 3265 1903
rect 3282 1856 3285 1966
rect 3294 1946 3297 2033
rect 3306 1983 3309 2156
rect 3314 2146 3317 2163
rect 3322 2153 3325 2206
rect 3330 2183 3333 2206
rect 3314 2143 3325 2146
rect 3322 2133 3325 2143
rect 3314 2013 3317 2126
rect 3330 2123 3333 2176
rect 3338 2153 3341 2313
rect 3370 2306 3373 2353
rect 3378 2313 3381 2416
rect 3394 2306 3397 2423
rect 3358 2303 3373 2306
rect 3386 2303 3397 2306
rect 3338 2106 3341 2136
rect 3346 2123 3349 2296
rect 3358 2246 3361 2303
rect 3354 2243 3361 2246
rect 3354 2223 3357 2243
rect 3354 2203 3357 2216
rect 3362 2203 3365 2226
rect 3354 2193 3365 2196
rect 3354 2133 3357 2146
rect 3362 2123 3365 2176
rect 3334 2103 3341 2106
rect 3258 1793 3265 1796
rect 3274 1853 3285 1856
rect 3290 1943 3297 1946
rect 3258 1736 3261 1793
rect 3274 1756 3277 1853
rect 3290 1813 3293 1943
rect 3314 1933 3317 1996
rect 3334 1956 3337 2103
rect 3346 2086 3349 2106
rect 3346 2083 3357 2086
rect 3354 2036 3357 2083
rect 3346 2033 3357 2036
rect 3334 1953 3341 1956
rect 3282 1793 3293 1796
rect 3298 1763 3301 1926
rect 3338 1923 3341 1953
rect 3346 1906 3349 2033
rect 3370 2006 3373 2286
rect 3386 2226 3389 2303
rect 3386 2223 3393 2226
rect 3378 2143 3381 2216
rect 3390 2176 3393 2223
rect 3386 2173 3393 2176
rect 3386 2126 3389 2173
rect 3382 2123 3389 2126
rect 3382 2056 3385 2123
rect 3382 2053 3389 2056
rect 3362 2003 3373 2006
rect 3342 1903 3349 1906
rect 3306 1813 3309 1826
rect 3314 1813 3317 1836
rect 3322 1806 3325 1816
rect 3306 1796 3309 1806
rect 3314 1803 3325 1806
rect 3306 1793 3317 1796
rect 3330 1793 3333 1826
rect 3342 1816 3345 1903
rect 3338 1813 3345 1816
rect 3274 1753 3301 1756
rect 3234 1653 3237 1726
rect 3242 1723 3245 1736
rect 3258 1733 3265 1736
rect 3234 1613 3237 1636
rect 3214 1493 3221 1496
rect 3174 1373 3181 1376
rect 3178 1356 3181 1373
rect 3178 1353 3189 1356
rect 3114 1113 3117 1146
rect 3162 1136 3165 1336
rect 3170 1333 3173 1346
rect 3170 1313 3173 1326
rect 3170 1143 3173 1306
rect 3186 1296 3189 1353
rect 3178 1293 3189 1296
rect 3114 1076 3117 1096
rect 3130 1083 3133 1126
rect 3114 1073 3121 1076
rect 3098 1023 3109 1026
rect 3098 833 3101 956
rect 3106 903 3109 1023
rect 3118 986 3121 1073
rect 3114 983 3121 986
rect 3114 933 3117 983
rect 3130 966 3133 1076
rect 3138 983 3141 1136
rect 3162 1133 3173 1136
rect 3146 1103 3149 1126
rect 3154 1123 3165 1126
rect 3170 1066 3173 1133
rect 3162 1063 3173 1066
rect 3122 963 3133 966
rect 3098 776 3101 816
rect 3106 803 3109 826
rect 3114 823 3117 836
rect 3082 773 3101 776
rect 3074 733 3077 756
rect 3082 723 3085 773
rect 3066 703 3077 706
rect 3074 616 3077 703
rect 3090 686 3093 756
rect 3098 693 3101 736
rect 3106 733 3109 796
rect 3114 726 3117 786
rect 3110 723 3117 726
rect 3090 683 3101 686
rect 3066 613 3077 616
rect 3050 603 3061 606
rect 3050 593 3053 603
rect 3066 596 3069 613
rect 3058 593 3069 596
rect 3042 583 3053 586
rect 3050 526 3053 583
rect 3058 533 3061 593
rect 3074 573 3077 596
rect 3066 533 3069 546
rect 3050 523 3077 526
rect 3074 506 3077 523
rect 3066 503 3077 506
rect 3066 436 3069 503
rect 3066 433 3077 436
rect 3042 413 3045 426
rect 3026 403 3037 406
rect 3026 336 3029 403
rect 3042 383 3045 406
rect 3066 403 3069 416
rect 3026 333 3037 336
rect 3018 296 3021 316
rect 3034 306 3037 333
rect 3042 313 3045 356
rect 3034 303 3045 306
rect 3018 293 3025 296
rect 3022 186 3025 293
rect 3034 203 3037 226
rect 3042 213 3045 303
rect 3050 283 3053 326
rect 3074 316 3077 433
rect 3082 333 3085 536
rect 3090 523 3093 546
rect 3098 473 3101 683
rect 3110 586 3113 723
rect 3122 603 3125 963
rect 3146 936 3149 1006
rect 3154 1003 3157 1016
rect 3130 933 3141 936
rect 3146 933 3157 936
rect 3130 823 3133 933
rect 3138 923 3149 926
rect 3138 803 3141 923
rect 3146 813 3149 856
rect 3154 813 3157 933
rect 3130 776 3133 796
rect 3130 773 3137 776
rect 3134 636 3137 773
rect 3130 633 3137 636
rect 3110 583 3117 586
rect 3114 466 3117 583
rect 3130 543 3133 633
rect 3138 533 3141 616
rect 3106 463 3117 466
rect 3098 423 3101 436
rect 3106 413 3109 463
rect 3122 413 3125 426
rect 3114 383 3117 406
rect 3050 203 3053 226
rect 3058 213 3061 236
rect 3022 183 3029 186
rect 3026 106 3029 183
rect 3066 136 3069 316
rect 3074 313 3085 316
rect 3082 166 3085 313
rect 3098 203 3101 326
rect 3106 303 3109 316
rect 3114 313 3117 336
rect 3106 213 3109 226
rect 3122 213 3125 396
rect 3138 346 3141 456
rect 3146 403 3149 806
rect 3154 726 3157 806
rect 3162 746 3165 1063
rect 3170 1003 3173 1056
rect 3170 793 3173 946
rect 3178 843 3181 1293
rect 3202 1276 3205 1326
rect 3194 1273 3205 1276
rect 3186 1196 3189 1226
rect 3194 1213 3197 1273
rect 3214 1246 3217 1493
rect 3226 1463 3229 1606
rect 3226 1403 3229 1416
rect 3226 1313 3229 1396
rect 3226 1253 3229 1276
rect 3214 1243 3221 1246
rect 3210 1216 3213 1226
rect 3202 1213 3213 1216
rect 3186 1193 3193 1196
rect 3190 1116 3193 1193
rect 3190 1113 3197 1116
rect 3186 933 3189 1106
rect 3194 943 3197 1113
rect 3202 1073 3205 1213
rect 3210 1143 3213 1206
rect 3218 1093 3221 1243
rect 3226 1213 3229 1246
rect 3234 1206 3237 1606
rect 3226 1203 3237 1206
rect 3226 1163 3229 1203
rect 3234 1133 3237 1196
rect 3242 1133 3245 1696
rect 3250 1613 3253 1726
rect 3262 1656 3265 1733
rect 3258 1653 3265 1656
rect 3258 1633 3261 1653
rect 3258 1526 3261 1616
rect 3266 1533 3269 1616
rect 3258 1523 3269 1526
rect 3274 1516 3277 1726
rect 3290 1606 3293 1686
rect 3298 1613 3301 1753
rect 3314 1746 3317 1793
rect 3314 1743 3321 1746
rect 3306 1633 3309 1736
rect 3318 1666 3321 1743
rect 3314 1663 3321 1666
rect 3314 1616 3317 1663
rect 3330 1646 3333 1726
rect 3310 1613 3317 1616
rect 3322 1643 3333 1646
rect 3290 1603 3301 1606
rect 3250 1423 3253 1516
rect 3266 1513 3277 1516
rect 3266 1426 3269 1513
rect 3282 1506 3285 1536
rect 3290 1523 3293 1536
rect 3298 1506 3301 1603
rect 3310 1546 3313 1613
rect 3310 1543 3317 1546
rect 3274 1503 3285 1506
rect 3294 1503 3301 1506
rect 3266 1423 3273 1426
rect 3250 1223 3253 1406
rect 3258 1353 3261 1416
rect 3270 1346 3273 1423
rect 3266 1343 3273 1346
rect 3282 1343 3285 1416
rect 3294 1386 3297 1503
rect 3294 1383 3301 1386
rect 3258 1213 3261 1336
rect 3266 1196 3269 1343
rect 3290 1336 3293 1366
rect 3282 1333 3293 1336
rect 3298 1333 3301 1383
rect 3274 1313 3277 1326
rect 3282 1223 3285 1333
rect 3274 1213 3293 1216
rect 3250 1193 3269 1196
rect 3250 1133 3253 1193
rect 3242 1086 3245 1126
rect 3210 1083 3245 1086
rect 3250 1123 3261 1126
rect 3202 973 3205 1036
rect 3210 1003 3213 1083
rect 3194 923 3197 936
rect 3186 913 3205 916
rect 3186 803 3189 906
rect 3194 783 3197 816
rect 3162 743 3181 746
rect 3194 733 3197 746
rect 3154 723 3165 726
rect 3154 703 3157 716
rect 3162 626 3165 723
rect 3186 643 3189 726
rect 3202 636 3205 886
rect 3210 803 3213 906
rect 3218 893 3221 1046
rect 3226 1003 3229 1016
rect 3242 986 3245 1006
rect 3238 983 3245 986
rect 3218 813 3221 836
rect 3154 623 3165 626
rect 3194 633 3205 636
rect 3154 593 3157 623
rect 3154 403 3157 546
rect 3138 343 3149 346
rect 3114 193 3117 206
rect 3130 203 3133 336
rect 3146 196 3149 343
rect 3162 303 3165 616
rect 3170 603 3189 606
rect 3194 573 3197 633
rect 3218 566 3221 736
rect 3226 723 3229 936
rect 3238 906 3241 983
rect 3250 953 3253 1123
rect 3266 1053 3269 1176
rect 3274 1136 3277 1206
rect 3282 1163 3285 1206
rect 3290 1153 3293 1213
rect 3274 1133 3285 1136
rect 3282 1046 3285 1133
rect 3298 1123 3301 1326
rect 3306 1323 3309 1526
rect 3314 1333 3317 1543
rect 3322 1526 3325 1643
rect 3338 1636 3341 1813
rect 3346 1783 3349 1806
rect 3354 1733 3357 1906
rect 3346 1713 3349 1726
rect 3330 1633 3341 1636
rect 3330 1533 3333 1633
rect 3338 1543 3341 1626
rect 3346 1603 3349 1616
rect 3346 1533 3349 1556
rect 3322 1523 3349 1526
rect 3322 1423 3325 1516
rect 3330 1513 3341 1516
rect 3346 1506 3349 1523
rect 3338 1503 3349 1506
rect 3338 1413 3341 1503
rect 3354 1496 3357 1616
rect 3350 1493 3357 1496
rect 3350 1436 3353 1493
rect 3346 1433 3353 1436
rect 3274 1043 3285 1046
rect 3250 913 3253 936
rect 3258 923 3261 1016
rect 3274 946 3277 1043
rect 3298 1023 3301 1036
rect 3282 1013 3301 1016
rect 3298 993 3301 1006
rect 3274 943 3281 946
rect 3238 903 3245 906
rect 3266 903 3269 936
rect 3234 706 3237 876
rect 3242 786 3245 903
rect 3278 896 3281 943
rect 3306 926 3309 1236
rect 3314 1203 3317 1276
rect 3322 1243 3325 1316
rect 3330 1273 3333 1336
rect 3314 1003 3317 1156
rect 3322 1133 3325 1226
rect 3322 1086 3325 1126
rect 3330 1106 3333 1256
rect 3338 1223 3341 1406
rect 3346 1396 3349 1433
rect 3354 1403 3357 1416
rect 3346 1393 3357 1396
rect 3346 1333 3349 1386
rect 3346 1233 3349 1326
rect 3354 1323 3357 1393
rect 3362 1306 3365 2003
rect 3370 1703 3373 1856
rect 3358 1303 3365 1306
rect 3358 1226 3361 1303
rect 3346 1223 3361 1226
rect 3338 1143 3341 1216
rect 3346 1173 3349 1223
rect 3354 1166 3357 1216
rect 3362 1193 3365 1204
rect 3370 1203 3373 1646
rect 3378 1503 3381 2036
rect 3378 1423 3381 1496
rect 3378 1323 3381 1406
rect 3378 1193 3381 1316
rect 3346 1163 3357 1166
rect 3362 1183 3381 1186
rect 3346 1136 3349 1163
rect 3338 1133 3349 1136
rect 3354 1133 3357 1146
rect 3338 1113 3341 1126
rect 3330 1103 3345 1106
rect 3322 1083 3333 1086
rect 3330 1006 3333 1083
rect 3322 1003 3333 1006
rect 3342 1006 3345 1103
rect 3342 1003 3349 1006
rect 3290 913 3293 926
rect 3306 923 3313 926
rect 3250 803 3253 816
rect 3242 783 3249 786
rect 3230 703 3237 706
rect 3230 636 3233 703
rect 3246 696 3249 783
rect 3226 633 3233 636
rect 3242 693 3249 696
rect 3226 596 3229 633
rect 3234 613 3237 626
rect 3226 593 3233 596
rect 3186 563 3221 566
rect 3170 333 3173 526
rect 3178 413 3181 426
rect 3170 303 3173 316
rect 3178 276 3181 316
rect 3138 193 3149 196
rect 3170 273 3181 276
rect 3138 173 3141 193
rect 3058 133 3069 136
rect 3074 163 3085 166
rect 3074 133 3077 163
rect 3098 123 3101 136
rect 3170 123 3173 273
rect 3186 266 3189 563
rect 3202 446 3205 536
rect 3218 533 3221 546
rect 3230 536 3233 593
rect 3230 533 3237 536
rect 3210 523 3221 526
rect 3226 453 3229 526
rect 3234 506 3237 533
rect 3242 523 3245 693
rect 3250 603 3253 616
rect 3234 503 3245 506
rect 3258 503 3261 896
rect 3274 893 3281 896
rect 3266 763 3269 806
rect 3274 786 3277 893
rect 3282 803 3285 816
rect 3290 803 3293 816
rect 3274 783 3281 786
rect 3266 623 3269 726
rect 3278 696 3281 783
rect 3290 733 3293 796
rect 3298 753 3301 916
rect 3310 836 3313 923
rect 3306 833 3313 836
rect 3298 703 3301 726
rect 3306 706 3309 833
rect 3314 723 3317 816
rect 3322 783 3325 1003
rect 3330 933 3333 946
rect 3306 703 3321 706
rect 3278 693 3301 696
rect 3298 636 3301 693
rect 3318 646 3321 703
rect 3318 643 3325 646
rect 3298 633 3309 636
rect 3266 556 3269 616
rect 3290 556 3293 616
rect 3306 613 3309 633
rect 3314 573 3317 626
rect 3322 586 3325 643
rect 3330 623 3333 926
rect 3338 793 3341 986
rect 3346 776 3349 1003
rect 3354 933 3357 1126
rect 3362 983 3365 1183
rect 3370 976 3373 1166
rect 3362 973 3373 976
rect 3354 903 3357 926
rect 3362 906 3365 973
rect 3370 913 3373 926
rect 3362 903 3369 906
rect 3366 846 3369 903
rect 3366 843 3373 846
rect 3342 773 3349 776
rect 3342 646 3345 773
rect 3342 643 3349 646
rect 3338 613 3341 626
rect 3346 606 3349 643
rect 3330 603 3349 606
rect 3346 586 3349 603
rect 3322 583 3333 586
rect 3266 553 3293 556
rect 3266 526 3269 553
rect 3274 533 3301 536
rect 3306 533 3309 556
rect 3266 523 3277 526
rect 3242 446 3245 503
rect 3194 413 3197 446
rect 3202 443 3221 446
rect 3210 413 3213 436
rect 3194 313 3197 336
rect 3202 323 3205 406
rect 3210 306 3213 406
rect 3218 396 3221 443
rect 3226 443 3245 446
rect 3226 413 3229 443
rect 3274 423 3277 523
rect 3290 513 3293 526
rect 3290 486 3293 506
rect 3286 483 3293 486
rect 3218 393 3225 396
rect 3178 263 3189 266
rect 3206 303 3213 306
rect 3178 133 3181 263
rect 3206 236 3209 303
rect 3222 296 3225 393
rect 3218 293 3225 296
rect 3206 233 3213 236
rect 3186 213 3197 216
rect 3194 203 3197 213
rect 3202 173 3205 216
rect 3210 213 3213 233
rect 3178 123 3189 126
rect 3218 123 3221 293
rect 3234 236 3237 416
rect 3242 413 3261 416
rect 3242 313 3245 413
rect 3250 366 3253 406
rect 3258 403 3261 413
rect 3274 366 3277 416
rect 3250 363 3277 366
rect 3258 333 3261 363
rect 3286 346 3289 483
rect 3286 343 3293 346
rect 3250 303 3253 316
rect 3266 286 3269 326
rect 3266 283 3277 286
rect 3226 233 3237 236
rect 3226 203 3229 233
rect 3250 203 3253 226
rect 3266 203 3269 226
rect 3274 203 3277 283
rect 3282 213 3285 326
rect 3290 306 3293 343
rect 3298 323 3301 533
rect 3330 526 3333 583
rect 3314 436 3317 526
rect 3322 523 3333 526
rect 3342 583 3349 586
rect 3354 586 3357 826
rect 3362 813 3365 826
rect 3362 783 3365 806
rect 3370 766 3373 843
rect 3366 763 3373 766
rect 3366 636 3369 763
rect 3366 633 3373 636
rect 3362 596 3365 616
rect 3370 603 3373 633
rect 3378 596 3381 1176
rect 3386 786 3389 2053
rect 3394 1773 3397 2156
rect 3394 1713 3397 1726
rect 3394 1643 3397 1706
rect 3394 1623 3397 1636
rect 3394 1533 3397 1546
rect 3394 1513 3397 1526
rect 3394 1373 3397 1506
rect 3394 1353 3397 1366
rect 3394 1013 3397 1346
rect 3394 803 3397 1006
rect 3402 863 3405 2276
rect 3386 783 3393 786
rect 3390 636 3393 783
rect 3362 593 3381 596
rect 3386 633 3393 636
rect 3354 583 3365 586
rect 3322 503 3325 523
rect 3342 456 3345 583
rect 3354 473 3357 576
rect 3362 466 3365 583
rect 3378 493 3381 516
rect 3386 483 3389 633
rect 3354 463 3365 466
rect 3342 453 3349 456
rect 3314 433 3341 436
rect 3306 396 3309 426
rect 3314 403 3317 433
rect 3330 396 3333 426
rect 3306 393 3333 396
rect 3314 326 3317 386
rect 3338 353 3341 426
rect 3346 396 3349 453
rect 3354 413 3357 463
rect 3370 446 3373 476
rect 3394 466 3397 616
rect 3366 443 3373 446
rect 3390 463 3397 466
rect 3346 393 3357 396
rect 3314 323 3333 326
rect 3290 303 3301 306
rect 3322 303 3325 316
rect 3298 226 3301 303
rect 3290 223 3301 226
rect 3290 206 3293 223
rect 3314 213 3317 226
rect 3330 213 3333 323
rect 3338 296 3341 346
rect 3354 326 3357 393
rect 3366 346 3369 443
rect 3366 343 3373 346
rect 3378 343 3381 426
rect 3354 323 3365 326
rect 3370 316 3373 343
rect 3390 336 3393 463
rect 3402 353 3405 826
rect 3390 333 3397 336
rect 3362 313 3373 316
rect 3338 293 3357 296
rect 3354 206 3357 293
rect 3378 213 3381 316
rect 3394 313 3397 333
rect 3282 203 3293 206
rect 3282 123 3285 203
rect 3322 196 3325 206
rect 3290 193 3325 196
rect 3338 203 3357 206
rect 3290 123 3293 193
rect 3298 133 3301 146
rect 3178 116 3181 123
rect 3162 113 3181 116
rect 3018 103 3029 106
rect 3306 103 3309 126
rect 3314 123 3317 136
rect 3338 123 3341 203
rect 2922 73 2933 76
rect 2930 43 2933 73
rect 3018 6 3021 103
rect 3414 37 3434 3303
rect 3438 13 3458 3327
rect 3010 3 3021 6
<< metal3 >>
rect 497 3272 1790 3277
rect 497 3252 502 3272
rect 169 3242 1462 3247
rect 2361 3232 2470 3237
rect 2361 3227 2366 3232
rect 433 3222 462 3227
rect 457 3217 462 3222
rect 521 3222 550 3227
rect 601 3222 718 3227
rect 985 3222 1014 3227
rect 521 3217 526 3222
rect 457 3212 526 3217
rect 1009 3217 1014 3222
rect 1073 3222 1102 3227
rect 2337 3222 2366 3227
rect 2465 3227 2470 3232
rect 2553 3232 2630 3237
rect 2681 3232 2798 3237
rect 2553 3227 2558 3232
rect 2465 3222 2558 3227
rect 2625 3227 2630 3232
rect 2625 3222 2718 3227
rect 1073 3217 1078 3222
rect 1009 3212 1078 3217
rect 2305 3212 2454 3217
rect 2585 3212 2614 3217
rect 2449 3207 2590 3212
rect 297 3202 342 3207
rect 625 3202 718 3207
rect 841 3202 934 3207
rect 841 3197 846 3202
rect 273 3192 398 3197
rect 817 3192 846 3197
rect 929 3197 934 3202
rect 1145 3202 1214 3207
rect 1273 3202 1374 3207
rect 2921 3202 3070 3207
rect 1145 3197 1150 3202
rect 929 3192 958 3197
rect 1121 3192 1150 3197
rect 1209 3197 1214 3202
rect 2921 3197 2926 3202
rect 1209 3192 1238 3197
rect 1417 3192 1510 3197
rect 1417 3187 1422 3192
rect 313 3182 342 3187
rect 337 3177 342 3182
rect 409 3182 1422 3187
rect 1505 3187 1510 3192
rect 1553 3192 1638 3197
rect 1993 3192 2118 3197
rect 2137 3192 2190 3197
rect 2201 3192 2318 3197
rect 2465 3192 2574 3197
rect 2649 3192 2742 3197
rect 2897 3192 2926 3197
rect 3065 3197 3070 3202
rect 3113 3202 3222 3207
rect 3113 3197 3118 3202
rect 3065 3192 3118 3197
rect 3217 3197 3222 3202
rect 3217 3192 3310 3197
rect 1553 3187 1558 3192
rect 1505 3182 1558 3187
rect 1633 3187 1638 3192
rect 2113 3187 2118 3192
rect 1633 3182 1982 3187
rect 2113 3182 2342 3187
rect 2737 3182 2974 3187
rect 409 3177 414 3182
rect 1977 3177 1982 3182
rect 2545 3177 2742 3182
rect 337 3172 414 3177
rect 1041 3172 1334 3177
rect 761 3167 894 3172
rect 1041 3167 1046 3172
rect 1329 3167 1334 3172
rect 1409 3172 1494 3177
rect 1409 3167 1414 3172
rect 673 3162 766 3167
rect 889 3162 1046 3167
rect 1057 3162 1270 3167
rect 1329 3162 1414 3167
rect 1489 3167 1494 3172
rect 1561 3172 1590 3177
rect 1977 3172 2102 3177
rect 1561 3167 1566 3172
rect 1489 3162 1566 3167
rect 1585 3167 1590 3172
rect 2097 3167 2102 3172
rect 2353 3172 2550 3177
rect 2817 3172 2886 3177
rect 2985 3172 3206 3177
rect 2353 3167 2358 3172
rect 2881 3167 2990 3172
rect 1585 3162 1806 3167
rect 2097 3162 2358 3167
rect 2561 3162 2862 3167
rect 3289 3162 3318 3167
rect 1057 3157 1062 3162
rect 777 3152 1062 3157
rect 1073 3152 1102 3157
rect 1209 3152 1254 3157
rect 1097 3147 1214 3152
rect 185 3142 254 3147
rect 441 3142 582 3147
rect 625 3142 790 3147
rect 865 3142 966 3147
rect 409 3132 478 3137
rect 577 3132 582 3142
rect 1233 3137 1238 3147
rect 801 3132 910 3137
rect 985 3132 1238 3137
rect 1265 3137 1270 3162
rect 2017 3152 2078 3157
rect 2377 3152 2542 3157
rect 2593 3152 2710 3157
rect 2825 3152 3158 3157
rect 3169 3152 3390 3157
rect 2705 3147 2830 3152
rect 1345 3142 1406 3147
rect 1449 3142 1494 3147
rect 1681 3142 1742 3147
rect 1913 3142 1982 3147
rect 2145 3142 2262 3147
rect 2361 3142 2686 3147
rect 2849 3142 2990 3147
rect 2001 3137 2102 3142
rect 2145 3137 2150 3142
rect 1265 3132 1382 3137
rect 1473 3132 2006 3137
rect 2097 3132 2150 3137
rect 2257 3137 2262 3142
rect 3033 3137 3102 3142
rect 2257 3132 2478 3137
rect 2521 3132 2614 3137
rect 2649 3132 2694 3137
rect 577 3127 782 3132
rect 1377 3127 1478 3132
rect 2713 3127 2718 3137
rect 2729 3132 2838 3137
rect 3001 3132 3038 3137
rect 3097 3132 3126 3137
rect 2833 3127 3006 3132
rect 777 3122 1046 3127
rect 1185 3122 1222 3127
rect 1809 3122 1974 3127
rect 1985 3122 2334 3127
rect 2449 3122 2718 3127
rect 3049 3122 3078 3127
rect 425 3112 918 3117
rect 953 3112 1006 3117
rect 1041 3107 1046 3122
rect 1241 3117 1358 3122
rect 1969 3117 1974 3122
rect 2329 3117 2454 3122
rect 3153 3117 3158 3152
rect 3249 3132 3358 3137
rect 1193 3112 1246 3117
rect 1353 3112 1382 3117
rect 1473 3112 1830 3117
rect 1969 3112 2206 3117
rect 2217 3112 2310 3117
rect 2481 3112 2614 3117
rect 2705 3112 2870 3117
rect 297 3102 406 3107
rect 777 3102 806 3107
rect 801 3097 806 3102
rect 881 3102 910 3107
rect 1041 3102 1222 3107
rect 1241 3102 1390 3107
rect 881 3097 886 3102
rect 801 3092 886 3097
rect 1217 3097 1222 3102
rect 1473 3097 1478 3112
rect 1825 3107 1830 3112
rect 2865 3107 2870 3112
rect 2953 3112 2982 3117
rect 3153 3112 3286 3117
rect 2953 3107 2958 3112
rect 1489 3102 1574 3107
rect 1825 3102 1958 3107
rect 1953 3097 1958 3102
rect 2065 3102 2094 3107
rect 2113 3102 2278 3107
rect 2385 3102 2430 3107
rect 2577 3102 2646 3107
rect 2865 3102 2958 3107
rect 2065 3097 2070 3102
rect 1217 3092 1246 3097
rect 1345 3092 1478 3097
rect 1489 3092 1526 3097
rect 1953 3092 2070 3097
rect 2321 3092 2494 3097
rect 3081 3092 3230 3097
rect 1241 3087 1350 3092
rect 441 3082 590 3087
rect 1593 3082 1774 3087
rect 1793 3082 1886 3087
rect 2105 3082 2246 3087
rect 2569 3082 2766 3087
rect 1489 3077 1598 3082
rect 1769 3077 1774 3082
rect 2289 3077 2494 3082
rect 865 3072 1022 3077
rect 865 3057 870 3072
rect 1017 3057 1022 3072
rect 1297 3072 1446 3077
rect 1465 3072 1494 3077
rect 1769 3072 1950 3077
rect 1969 3072 2086 3077
rect 2265 3072 2294 3077
rect 2489 3072 2518 3077
rect 3137 3072 3398 3077
rect 1297 3067 1302 3072
rect 1041 3062 1110 3067
rect 1145 3062 1214 3067
rect 1273 3062 1302 3067
rect 1441 3067 1446 3072
rect 1617 3067 1750 3072
rect 1969 3067 1974 3072
rect 1441 3062 1622 3067
rect 1745 3062 1974 3067
rect 2081 3067 2086 3072
rect 2081 3062 2590 3067
rect 1145 3057 1150 3062
rect 377 3052 454 3057
rect 537 3052 654 3057
rect 841 3052 870 3057
rect 921 3052 998 3057
rect 1017 3052 1150 3057
rect 1209 3057 1214 3062
rect 1321 3057 1422 3062
rect 1209 3052 1238 3057
rect 1265 3052 1326 3057
rect 1417 3052 1502 3057
rect 1569 3052 1998 3057
rect 2089 3052 2174 3057
rect 2257 3052 2446 3057
rect 2601 3052 2694 3057
rect 537 3047 542 3052
rect 249 3042 542 3047
rect 649 3047 654 3052
rect 921 3047 926 3052
rect 649 3042 678 3047
rect 809 3042 926 3047
rect 993 3047 998 3052
rect 993 3042 1078 3047
rect 1265 3037 1270 3052
rect 2257 3047 2262 3052
rect 2441 3047 2606 3052
rect 1289 3042 1790 3047
rect 1929 3042 2262 3047
rect 2273 3042 2422 3047
rect 3209 3042 3246 3047
rect 1785 3037 1934 3042
rect 313 3032 398 3037
rect 553 3032 702 3037
rect 937 3032 1270 3037
rect 1409 3032 1598 3037
rect 2169 3032 2334 3037
rect 2369 3032 2406 3037
rect 2473 3032 2662 3037
rect 3105 3032 3198 3037
rect 3257 3032 3286 3037
rect 801 3027 870 3032
rect 1625 3027 1734 3032
rect 2473 3027 2478 3032
rect 401 3022 454 3027
rect 617 3022 742 3027
rect 777 3022 806 3027
rect 865 3022 1094 3027
rect 1297 3022 1446 3027
rect 1609 3022 1630 3027
rect 1729 3022 1774 3027
rect 1809 3022 1926 3027
rect 2009 3022 2118 3027
rect 1441 3017 1446 3022
rect 1529 3017 1614 3022
rect 2009 3017 2014 3022
rect 473 3012 558 3017
rect 673 3012 854 3017
rect 929 3012 966 3017
rect 1113 3012 1278 3017
rect 1305 3012 1334 3017
rect 1369 3012 1422 3017
rect 1441 3012 1534 3017
rect 1641 3012 1782 3017
rect 1793 3012 2014 3017
rect 2113 3017 2118 3022
rect 2193 3022 2438 3027
rect 2449 3022 2478 3027
rect 2657 3027 2662 3032
rect 3193 3027 3262 3032
rect 2657 3022 2686 3027
rect 2865 3022 2950 3027
rect 2193 3017 2198 3022
rect 2433 3017 2438 3022
rect 2113 3012 2198 3017
rect 2209 3012 2318 3017
rect 2377 3012 2406 3017
rect 2433 3012 2678 3017
rect 2857 3012 2886 3017
rect 961 3007 1118 3012
rect 1273 3007 1278 3012
rect 2881 3007 2886 3012
rect 2953 3012 3126 3017
rect 3209 3012 3318 3017
rect 2953 3007 2958 3012
rect 3121 3007 3126 3012
rect 721 3002 950 3007
rect 1273 3002 1350 3007
rect 1553 3002 1694 3007
rect 1705 3002 1838 3007
rect 1857 3002 1878 3007
rect 2025 3002 2182 3007
rect 2265 3002 2374 3007
rect 2505 3002 2542 3007
rect 2881 3002 2958 3007
rect 2977 3002 3110 3007
rect 3121 3002 3278 3007
rect 3353 3002 3398 3007
rect 1665 2997 1670 3002
rect 1857 2997 1862 3002
rect 137 2992 222 2997
rect 305 2992 406 2997
rect 561 2992 630 2997
rect 681 2992 902 2997
rect 993 2992 1358 2997
rect 1393 2992 1510 2997
rect 1665 2992 1862 2997
rect 1889 2992 1926 2997
rect 1945 2992 2134 2997
rect 2177 2992 2286 2997
rect 1921 2987 1926 2992
rect 2177 2987 2182 2992
rect 2369 2987 2374 3002
rect 2393 2992 2494 2997
rect 2553 2992 2718 2997
rect 3097 2992 3222 2997
rect 209 2982 366 2987
rect 441 2982 518 2987
rect 593 2982 798 2987
rect 873 2982 926 2987
rect 961 2982 1406 2987
rect 1433 2982 1526 2987
rect 1577 2982 1902 2987
rect 1921 2982 2070 2987
rect 2121 2982 2182 2987
rect 2305 2982 2350 2987
rect 2369 2982 2566 2987
rect 3057 2982 3246 2987
rect 209 2977 214 2982
rect 193 2972 214 2977
rect 233 2972 262 2977
rect 497 2972 622 2977
rect 689 2972 830 2977
rect 889 2972 1038 2977
rect 1089 2972 1254 2977
rect 1329 2972 1358 2977
rect 257 2967 262 2972
rect 377 2967 502 2972
rect 1353 2967 1358 2972
rect 1425 2972 1734 2977
rect 1937 2972 2086 2977
rect 2289 2972 2622 2977
rect 2641 2972 2710 2977
rect 1425 2967 1430 2972
rect 1753 2967 1942 2972
rect 2641 2967 2646 2972
rect 257 2962 382 2967
rect 521 2962 574 2967
rect 657 2962 990 2967
rect 1161 2962 1278 2967
rect 1353 2962 1430 2967
rect 1449 2962 1558 2967
rect 1681 2962 1758 2967
rect 1961 2962 2358 2967
rect 2553 2962 2646 2967
rect 2705 2967 2710 2972
rect 2753 2972 2918 2977
rect 2753 2967 2758 2972
rect 2705 2962 2758 2967
rect 2913 2967 2918 2972
rect 2913 2962 3126 2967
rect 505 2952 574 2957
rect 633 2952 662 2957
rect 777 2952 838 2957
rect 865 2952 894 2957
rect 1009 2952 1158 2957
rect 1233 2952 1302 2957
rect 1513 2952 2206 2957
rect 2345 2952 2470 2957
rect 2521 2952 2694 2957
rect 657 2947 782 2952
rect 129 2942 246 2947
rect 273 2942 430 2947
rect 257 2932 286 2937
rect 281 2917 286 2932
rect 441 2932 518 2937
rect 713 2932 774 2937
rect 441 2917 446 2932
rect 801 2927 806 2952
rect 825 2942 854 2947
rect 1137 2942 1430 2947
rect 1441 2942 1502 2947
rect 1569 2942 1942 2947
rect 1961 2942 2054 2947
rect 2129 2942 2310 2947
rect 2441 2942 2614 2947
rect 849 2937 1030 2942
rect 1497 2937 1574 2942
rect 1937 2937 1942 2942
rect 1025 2932 1102 2937
rect 1153 2932 1182 2937
rect 1225 2932 1342 2937
rect 1593 2932 1894 2937
rect 1937 2932 1990 2937
rect 2065 2932 2270 2937
rect 2321 2932 2366 2937
rect 2481 2932 2686 2937
rect 521 2922 702 2927
rect 801 2922 1014 2927
rect 1201 2922 1278 2927
rect 1313 2922 1582 2927
rect 1825 2922 1974 2927
rect 1993 2922 2054 2927
rect 281 2912 446 2917
rect 697 2917 702 2922
rect 1033 2917 1126 2922
rect 1577 2917 1830 2922
rect 2065 2917 2070 2932
rect 2769 2927 2774 2947
rect 2801 2942 2902 2947
rect 3201 2942 3238 2947
rect 2921 2937 2990 2942
rect 2881 2932 2926 2937
rect 2985 2932 3222 2937
rect 3241 2932 3262 2937
rect 2217 2922 2278 2927
rect 2457 2922 2550 2927
rect 2665 2922 2870 2927
rect 697 2912 886 2917
rect 897 2912 950 2917
rect 961 2912 1038 2917
rect 1121 2912 1150 2917
rect 1161 2912 1398 2917
rect 1849 2912 1878 2917
rect 897 2907 902 2912
rect 1873 2907 1878 2912
rect 1953 2912 2070 2917
rect 2201 2912 2230 2917
rect 2361 2912 2398 2917
rect 2545 2912 2550 2922
rect 2865 2917 2870 2922
rect 2945 2922 2974 2927
rect 2945 2917 2950 2922
rect 2721 2912 2758 2917
rect 2865 2912 2950 2917
rect 3217 2912 3286 2917
rect 1953 2907 1958 2912
rect 465 2902 630 2907
rect 841 2902 902 2907
rect 969 2902 1262 2907
rect 1273 2902 1326 2907
rect 1361 2902 1550 2907
rect 1545 2897 1550 2902
rect 1633 2902 1662 2907
rect 1705 2902 1846 2907
rect 1873 2902 1958 2907
rect 1977 2902 2006 2907
rect 1633 2897 1638 2902
rect 489 2892 526 2897
rect 521 2887 526 2892
rect 625 2892 742 2897
rect 777 2892 1030 2897
rect 625 2887 630 2892
rect 1025 2887 1030 2892
rect 1153 2892 1206 2897
rect 1281 2892 1470 2897
rect 1545 2892 1638 2897
rect 2001 2897 2006 2902
rect 2081 2902 2238 2907
rect 2313 2902 2390 2907
rect 2505 2902 2606 2907
rect 3025 2902 3262 2907
rect 2081 2897 2086 2902
rect 2001 2892 2086 2897
rect 2177 2892 2286 2897
rect 2353 2892 2494 2897
rect 2601 2892 2630 2897
rect 2745 2892 3166 2897
rect 1153 2887 1158 2892
rect 2489 2887 2606 2892
rect 3161 2887 3166 2892
rect 3289 2892 3318 2897
rect 3289 2887 3294 2892
rect 521 2882 630 2887
rect 913 2882 1006 2887
rect 1025 2882 1158 2887
rect 1177 2882 1390 2887
rect 1657 2882 1790 2887
rect 2241 2882 2398 2887
rect 3089 2882 3142 2887
rect 3161 2882 3294 2887
rect 361 2872 502 2877
rect 649 2872 798 2877
rect 841 2872 862 2877
rect 1329 2872 1502 2877
rect 2049 2872 2158 2877
rect 649 2867 654 2872
rect 625 2862 654 2867
rect 793 2867 798 2872
rect 1129 2867 1310 2872
rect 2049 2867 2054 2872
rect 793 2862 886 2867
rect 1073 2862 1134 2867
rect 1305 2862 1598 2867
rect 1929 2862 2054 2867
rect 2153 2867 2158 2872
rect 2353 2872 2502 2877
rect 2153 2862 2230 2867
rect 2225 2857 2230 2862
rect 2353 2857 2358 2872
rect 2497 2867 2502 2872
rect 2601 2872 2854 2877
rect 3049 2872 3078 2877
rect 2601 2867 2606 2872
rect 2377 2862 2438 2867
rect 2497 2862 2606 2867
rect 481 2852 534 2857
rect 617 2852 662 2857
rect 705 2852 926 2857
rect 1145 2852 1678 2857
rect 1697 2852 1902 2857
rect 2225 2852 2358 2857
rect 2433 2857 2438 2862
rect 2433 2852 2478 2857
rect 2873 2852 3006 2857
rect 1697 2847 1702 2852
rect 609 2842 678 2847
rect 961 2842 1054 2847
rect 1185 2842 1254 2847
rect 1377 2842 1406 2847
rect 1649 2842 1702 2847
rect 1897 2847 1902 2852
rect 1897 2842 2174 2847
rect 2625 2842 2838 2847
rect 825 2837 918 2842
rect 961 2837 966 2842
rect 337 2832 406 2837
rect 337 2827 342 2832
rect 185 2822 342 2827
rect 401 2827 406 2832
rect 529 2832 566 2837
rect 665 2832 702 2837
rect 713 2832 830 2837
rect 913 2832 966 2837
rect 1049 2837 1054 2842
rect 1401 2837 1654 2842
rect 1769 2837 1862 2842
rect 2873 2837 2878 2852
rect 1049 2832 1214 2837
rect 1673 2832 1726 2837
rect 1745 2832 1774 2837
rect 1857 2832 1886 2837
rect 2417 2832 2446 2837
rect 2825 2832 2878 2837
rect 3001 2837 3006 2852
rect 3049 2842 3206 2847
rect 3049 2837 3054 2842
rect 3001 2832 3054 2837
rect 3201 2837 3206 2842
rect 3201 2832 3230 2837
rect 529 2827 534 2832
rect 401 2822 534 2827
rect 553 2822 582 2827
rect 649 2822 878 2827
rect 985 2822 1086 2827
rect 1321 2822 1430 2827
rect 1449 2822 1550 2827
rect 1105 2817 1278 2822
rect 1321 2817 1326 2822
rect 89 2812 206 2817
rect 353 2812 382 2817
rect 529 2812 870 2817
rect 881 2812 950 2817
rect 1001 2812 1110 2817
rect 1273 2812 1326 2817
rect 1425 2817 1430 2822
rect 1593 2817 1686 2822
rect 1425 2812 1598 2817
rect 1681 2812 1710 2817
rect 377 2807 534 2812
rect 1745 2807 1750 2832
rect 3073 2827 3174 2832
rect 1769 2822 1878 2827
rect 1905 2822 2134 2827
rect 1905 2817 1910 2822
rect 1793 2812 1910 2817
rect 2129 2817 2134 2822
rect 2193 2822 2398 2827
rect 2193 2817 2198 2822
rect 2129 2812 2198 2817
rect 2393 2817 2398 2822
rect 2465 2822 2534 2827
rect 2633 2822 2742 2827
rect 2817 2822 2950 2827
rect 2993 2822 3078 2827
rect 3169 2822 3198 2827
rect 2465 2817 2470 2822
rect 2393 2812 2470 2817
rect 2529 2817 2534 2822
rect 2529 2812 2558 2817
rect 2977 2812 3070 2817
rect 3105 2812 3214 2817
rect 1929 2807 2094 2812
rect 553 2802 774 2807
rect 929 2802 1750 2807
rect 1897 2802 1934 2807
rect 2089 2802 2118 2807
rect 2697 2802 2798 2807
rect 3177 2802 3238 2807
rect 3305 2802 3382 2807
rect 769 2797 934 2802
rect 121 2792 438 2797
rect 481 2792 750 2797
rect 953 2792 1094 2797
rect 1329 2792 1510 2797
rect 1585 2792 1894 2797
rect 1905 2792 1926 2797
rect 1969 2792 2790 2797
rect 1201 2787 1302 2792
rect 329 2782 382 2787
rect 417 2782 550 2787
rect 569 2782 1206 2787
rect 1297 2782 1390 2787
rect 1633 2782 1950 2787
rect 545 2772 550 2782
rect 1969 2777 2078 2782
rect 2233 2777 2302 2782
rect 689 2772 846 2777
rect 945 2772 1030 2777
rect 1217 2772 1270 2777
rect 545 2767 670 2772
rect 1025 2767 1222 2772
rect 1265 2767 1270 2772
rect 1337 2772 1446 2777
rect 1457 2772 1782 2777
rect 1921 2772 1974 2777
rect 2073 2772 2238 2777
rect 2297 2772 2326 2777
rect 2337 2772 2382 2777
rect 2457 2772 2606 2777
rect 2849 2772 3038 2777
rect 1337 2767 1342 2772
rect 121 2762 254 2767
rect 665 2762 702 2767
rect 873 2762 1006 2767
rect 1265 2762 1342 2767
rect 1441 2767 1446 2772
rect 1441 2762 1470 2767
rect 1625 2762 1710 2767
rect 1865 2762 2062 2767
rect 2249 2762 2278 2767
rect 121 2757 126 2762
rect 89 2752 126 2757
rect 249 2757 254 2762
rect 1465 2757 1558 2762
rect 2057 2757 2254 2762
rect 2321 2757 2326 2772
rect 2849 2757 2854 2772
rect 249 2752 310 2757
rect 609 2752 814 2757
rect 985 2752 1062 2757
rect 1137 2752 1230 2757
rect 1553 2752 2038 2757
rect 2321 2752 2854 2757
rect 3033 2757 3038 2772
rect 3033 2752 3062 2757
rect 2033 2747 2038 2752
rect 137 2742 246 2747
rect 425 2742 478 2747
rect 617 2742 838 2747
rect 913 2742 998 2747
rect 1009 2742 1094 2747
rect 1185 2742 1542 2747
rect 1665 2742 1694 2747
rect 1721 2742 1830 2747
rect 1897 2742 1974 2747
rect 2033 2742 2118 2747
rect 2161 2742 2310 2747
rect 2505 2742 2558 2747
rect 689 2737 694 2742
rect 1009 2737 1014 2742
rect 1185 2737 1190 2742
rect 1537 2737 1670 2742
rect 2113 2737 2118 2742
rect 2305 2737 2438 2742
rect 2505 2737 2510 2742
rect 353 2732 422 2737
rect 457 2732 526 2737
rect 665 2732 694 2737
rect 761 2732 886 2737
rect 905 2732 1014 2737
rect 1049 2732 1150 2737
rect 1161 2732 1190 2737
rect 1809 2732 1862 2737
rect 2113 2732 2182 2737
rect 2433 2732 2510 2737
rect 2553 2737 2558 2742
rect 2625 2742 2654 2747
rect 2865 2742 3166 2747
rect 2625 2737 2630 2742
rect 2553 2732 2630 2737
rect 545 2727 646 2732
rect 881 2727 886 2732
rect 1697 2727 1774 2732
rect 1881 2727 2014 2732
rect 457 2722 550 2727
rect 641 2722 678 2727
rect 881 2722 958 2727
rect 1025 2722 1134 2727
rect 1177 2722 1270 2727
rect 1345 2722 1486 2727
rect 1513 2722 1702 2727
rect 1769 2722 1886 2727
rect 2009 2722 2198 2727
rect 2369 2722 2414 2727
rect 3289 2722 3350 2727
rect 1025 2717 1030 2722
rect 249 2712 398 2717
rect 537 2712 638 2717
rect 753 2712 838 2717
rect 849 2712 1030 2717
rect 1041 2712 1102 2717
rect 1249 2712 1318 2717
rect 1385 2712 1414 2717
rect 833 2707 838 2712
rect 489 2702 558 2707
rect 601 2702 662 2707
rect 833 2702 862 2707
rect 889 2702 1014 2707
rect 281 2697 382 2702
rect 1009 2697 1014 2702
rect 1113 2702 1174 2707
rect 1113 2697 1118 2702
rect 257 2692 286 2697
rect 377 2692 406 2697
rect 433 2692 566 2697
rect 825 2692 982 2697
rect 1009 2692 1118 2697
rect 1409 2697 1414 2712
rect 1713 2712 1758 2717
rect 1841 2712 2150 2717
rect 2209 2712 2350 2717
rect 2545 2712 2638 2717
rect 2817 2712 2958 2717
rect 3017 2712 3150 2717
rect 1713 2697 1718 2712
rect 2145 2707 2214 2712
rect 1737 2702 2126 2707
rect 2329 2702 2414 2707
rect 2721 2702 2838 2707
rect 3313 2702 3398 2707
rect 1409 2692 1718 2697
rect 1961 2692 1990 2697
rect 2137 2692 2318 2697
rect 2657 2692 2686 2697
rect 2897 2692 3078 2697
rect 1985 2687 2142 2692
rect 2681 2687 2766 2692
rect 2897 2687 2902 2692
rect 233 2682 534 2687
rect 1873 2682 1950 2687
rect 849 2677 950 2682
rect 1945 2677 1950 2682
rect 2185 2682 2214 2687
rect 2433 2682 2542 2687
rect 2761 2682 2902 2687
rect 3073 2687 3078 2692
rect 3161 2692 3214 2697
rect 3281 2692 3366 2697
rect 3161 2687 3166 2692
rect 3073 2682 3166 2687
rect 2185 2677 2190 2682
rect 2433 2677 2438 2682
rect 825 2672 854 2677
rect 945 2672 1198 2677
rect 1881 2672 1910 2677
rect 1945 2672 2190 2677
rect 2225 2672 2438 2677
rect 2537 2677 2542 2682
rect 2537 2672 2614 2677
rect 2649 2672 2742 2677
rect 265 2667 454 2672
rect 241 2662 270 2667
rect 449 2662 478 2667
rect 529 2662 630 2667
rect 689 2662 790 2667
rect 833 2662 934 2667
rect 529 2657 534 2662
rect 689 2657 694 2662
rect 1905 2657 1910 2672
rect 2225 2657 2230 2672
rect 2937 2662 2998 2667
rect 2329 2657 2406 2662
rect 249 2652 534 2657
rect 545 2652 694 2657
rect 705 2652 1046 2657
rect 1905 2652 2230 2657
rect 2305 2652 2334 2657
rect 2401 2652 2526 2657
rect 705 2647 710 2652
rect 129 2642 238 2647
rect 377 2642 710 2647
rect 721 2642 806 2647
rect 921 2642 966 2647
rect 1057 2642 1310 2647
rect 2361 2642 2390 2647
rect 233 2637 238 2642
rect 297 2637 382 2642
rect 721 2637 726 2642
rect 961 2637 1062 2642
rect 2385 2637 2390 2642
rect 2537 2642 2694 2647
rect 2889 2642 2958 2647
rect 3009 2642 3118 2647
rect 2537 2637 2542 2642
rect 233 2632 302 2637
rect 401 2632 574 2637
rect 665 2632 726 2637
rect 745 2632 846 2637
rect 913 2632 942 2637
rect 2177 2632 2302 2637
rect 2385 2632 2542 2637
rect 2737 2632 2966 2637
rect 3217 2632 3278 2637
rect 2177 2627 2182 2632
rect 129 2622 182 2627
rect 321 2622 398 2627
rect 465 2622 558 2627
rect 793 2622 838 2627
rect 849 2622 1030 2627
rect 1105 2622 1142 2627
rect 1609 2622 1662 2627
rect 1721 2622 1822 2627
rect 1841 2622 2006 2627
rect 2057 2622 2182 2627
rect 2297 2627 2302 2632
rect 2297 2622 2326 2627
rect 2745 2622 2822 2627
rect 2873 2622 2982 2627
rect 273 2612 422 2617
rect 601 2612 670 2617
rect 713 2612 1014 2617
rect 1025 2612 1030 2622
rect 1721 2617 1726 2622
rect 1361 2612 1478 2617
rect 1697 2612 1726 2617
rect 1817 2617 1822 2622
rect 1817 2612 1862 2617
rect 2193 2612 2558 2617
rect 2657 2612 2686 2617
rect 2849 2612 2878 2617
rect 2961 2612 2990 2617
rect 201 2602 262 2607
rect 569 2602 590 2607
rect 625 2602 694 2607
rect 777 2602 822 2607
rect 905 2602 958 2607
rect 1161 2602 1246 2607
rect 1497 2602 1590 2607
rect 1977 2602 2206 2607
rect 2329 2602 2422 2607
rect 257 2597 262 2602
rect 1161 2597 1166 2602
rect 129 2592 222 2597
rect 257 2592 518 2597
rect 633 2592 894 2597
rect 969 2592 1078 2597
rect 1089 2592 1166 2597
rect 1241 2597 1246 2602
rect 1305 2597 1502 2602
rect 1585 2597 1590 2602
rect 1737 2597 1822 2602
rect 2201 2597 2334 2602
rect 1241 2592 1270 2597
rect 1281 2592 1310 2597
rect 1585 2592 1662 2597
rect 1713 2592 1742 2597
rect 1817 2592 1886 2597
rect 2153 2592 2182 2597
rect 889 2587 974 2592
rect 2177 2587 2182 2592
rect 2353 2592 2382 2597
rect 2353 2587 2358 2592
rect 489 2582 606 2587
rect 641 2582 862 2587
rect 1025 2582 1806 2587
rect 1801 2577 1806 2582
rect 1897 2582 2014 2587
rect 2057 2582 2150 2587
rect 2177 2582 2358 2587
rect 2657 2582 2662 2612
rect 2873 2607 2966 2612
rect 2705 2602 2774 2607
rect 3273 2602 3342 2607
rect 3273 2597 3278 2602
rect 2713 2592 2790 2597
rect 2881 2592 2966 2597
rect 2977 2592 3046 2597
rect 3177 2592 3214 2597
rect 3249 2592 3278 2597
rect 3337 2597 3342 2602
rect 3337 2592 3366 2597
rect 3273 2582 3310 2587
rect 1897 2577 1902 2582
rect 193 2572 286 2577
rect 529 2572 558 2577
rect 665 2572 902 2577
rect 913 2572 942 2577
rect 993 2572 1126 2577
rect 1145 2572 1206 2577
rect 1257 2572 1470 2577
rect 1497 2572 1718 2577
rect 1801 2572 1902 2577
rect 2929 2572 3078 2577
rect 3297 2572 3334 2577
rect 553 2567 670 2572
rect 913 2567 918 2572
rect 1441 2567 1446 2572
rect 441 2562 510 2567
rect 441 2557 446 2562
rect 417 2552 446 2557
rect 505 2557 510 2562
rect 753 2562 918 2567
rect 929 2562 1222 2567
rect 1441 2562 1694 2567
rect 2801 2562 2886 2567
rect 753 2557 758 2562
rect 1241 2557 1422 2562
rect 2801 2557 2806 2562
rect 505 2552 566 2557
rect 601 2552 758 2557
rect 777 2552 974 2557
rect 1105 2552 1246 2557
rect 1417 2552 1518 2557
rect 1649 2552 1678 2557
rect 2113 2552 2270 2557
rect 2777 2552 2806 2557
rect 2881 2557 2886 2562
rect 2929 2557 2934 2572
rect 2881 2552 2934 2557
rect 3073 2557 3078 2572
rect 3097 2562 3142 2567
rect 3241 2562 3326 2567
rect 3073 2552 3286 2557
rect 3329 2552 3390 2557
rect 89 2542 422 2547
rect 465 2542 502 2547
rect 601 2542 718 2547
rect 833 2542 934 2547
rect 1057 2542 1422 2547
rect 1529 2542 1598 2547
rect 1617 2537 1622 2547
rect 577 2532 638 2537
rect 1065 2532 1294 2537
rect 1393 2532 1510 2537
rect 1569 2532 1622 2537
rect 1649 2537 1654 2552
rect 1681 2542 1766 2547
rect 1857 2542 1966 2547
rect 2073 2542 2134 2547
rect 2601 2542 2678 2547
rect 2745 2542 3254 2547
rect 3265 2542 3382 2547
rect 1649 2532 1694 2537
rect 2089 2532 2118 2537
rect 465 2527 582 2532
rect 1617 2527 1622 2532
rect 2129 2527 2134 2542
rect 2497 2532 2846 2537
rect 2857 2532 2926 2537
rect 3049 2532 3158 2537
rect 193 2522 214 2527
rect 225 2522 470 2527
rect 593 2522 662 2527
rect 905 2522 1558 2527
rect 1617 2522 1790 2527
rect 1929 2522 2102 2527
rect 2129 2522 2302 2527
rect 2401 2522 2486 2527
rect 193 2497 198 2522
rect 2481 2517 2486 2522
rect 2617 2522 2654 2527
rect 2713 2522 3158 2527
rect 3177 2522 3246 2527
rect 2617 2517 2622 2522
rect 3241 2517 3246 2522
rect 3321 2522 3350 2527
rect 3321 2517 3326 2522
rect 257 2512 286 2517
rect 281 2497 286 2512
rect 481 2512 894 2517
rect 1033 2512 1150 2517
rect 1209 2512 1662 2517
rect 1753 2512 1822 2517
rect 2065 2512 2150 2517
rect 2481 2512 2622 2517
rect 2641 2512 3006 2517
rect 3041 2512 3118 2517
rect 481 2497 486 2512
rect 889 2507 1038 2512
rect 3113 2507 3118 2512
rect 3193 2512 3222 2517
rect 3241 2512 3326 2517
rect 3193 2507 3198 2512
rect 513 2502 670 2507
rect 1057 2502 1254 2507
rect 1313 2502 1414 2507
rect 1457 2502 1590 2507
rect 1649 2502 1742 2507
rect 1753 2502 2094 2507
rect 2649 2502 2678 2507
rect 1585 2497 1590 2502
rect 2673 2497 2678 2502
rect 2857 2502 2942 2507
rect 3113 2502 3198 2507
rect 3361 2502 3382 2507
rect 2857 2497 2862 2502
rect 193 2492 254 2497
rect 281 2492 486 2497
rect 505 2492 614 2497
rect 681 2492 1118 2497
rect 1225 2492 1478 2497
rect 1585 2492 1686 2497
rect 2073 2492 2118 2497
rect 2369 2492 2454 2497
rect 2673 2492 2862 2497
rect 3017 2492 3094 2497
rect 609 2487 686 2492
rect 561 2482 590 2487
rect 585 2477 590 2482
rect 761 2482 790 2487
rect 1009 2482 1134 2487
rect 1265 2482 1310 2487
rect 1473 2482 1502 2487
rect 1537 2482 1838 2487
rect 1905 2482 2166 2487
rect 2281 2482 2430 2487
rect 761 2477 766 2482
rect 1305 2477 1478 2482
rect 1905 2477 1910 2482
rect 585 2472 766 2477
rect 873 2472 1094 2477
rect 1169 2472 1286 2477
rect 1633 2472 1742 2477
rect 1737 2467 1742 2472
rect 1841 2472 1910 2477
rect 2169 2472 2366 2477
rect 1841 2467 1846 2472
rect 945 2462 990 2467
rect 1337 2462 1470 2467
rect 1609 2462 1662 2467
rect 1737 2462 1846 2467
rect 1865 2462 2054 2467
rect 2457 2462 2926 2467
rect 1081 2457 1318 2462
rect 977 2452 1086 2457
rect 1313 2452 1654 2457
rect 433 2442 966 2447
rect 1097 2442 1166 2447
rect 1209 2442 1302 2447
rect 1393 2442 1446 2447
rect 961 2437 1102 2442
rect 1649 2437 1654 2452
rect 2121 2452 2262 2457
rect 2121 2447 2126 2452
rect 1689 2442 1718 2447
rect 1921 2442 2126 2447
rect 2257 2447 2262 2452
rect 2457 2447 2462 2462
rect 2921 2457 2926 2462
rect 2921 2452 3070 2457
rect 3065 2447 3070 2452
rect 2257 2442 2286 2447
rect 2305 2442 2414 2447
rect 2433 2442 2462 2447
rect 2481 2442 2822 2447
rect 3065 2442 3390 2447
rect 2305 2437 2310 2442
rect 1121 2432 1238 2437
rect 1305 2432 1406 2437
rect 1649 2432 1862 2437
rect 2137 2432 2310 2437
rect 2409 2437 2414 2442
rect 2481 2437 2486 2442
rect 2409 2432 2486 2437
rect 2817 2437 2822 2442
rect 2817 2432 2910 2437
rect 2577 2427 2798 2432
rect 809 2422 958 2427
rect 1073 2422 1318 2427
rect 1417 2422 1550 2427
rect 1673 2422 1774 2427
rect 809 2417 814 2422
rect 337 2412 814 2417
rect 953 2417 958 2422
rect 1769 2417 1774 2422
rect 1857 2422 2086 2427
rect 2121 2422 2222 2427
rect 2233 2422 2358 2427
rect 2385 2422 2406 2427
rect 2441 2422 2582 2427
rect 2793 2422 2918 2427
rect 2937 2422 3054 2427
rect 1857 2417 1862 2422
rect 953 2412 982 2417
rect 1193 2412 1310 2417
rect 1353 2412 1478 2417
rect 1489 2412 1718 2417
rect 1769 2412 1862 2417
rect 2081 2417 2086 2422
rect 2401 2417 2406 2422
rect 2081 2412 2110 2417
rect 2217 2412 2246 2417
rect 2401 2412 2470 2417
rect 2593 2412 2830 2417
rect 2977 2412 3094 2417
rect 3305 2412 3350 2417
rect 1097 2407 1174 2412
rect 2105 2407 2222 2412
rect 2849 2407 2958 2412
rect 825 2402 1102 2407
rect 1169 2402 1222 2407
rect 1273 2402 1598 2407
rect 1617 2402 1678 2407
rect 1697 2402 1750 2407
rect 1881 2402 2014 2407
rect 2313 2402 2854 2407
rect 2953 2402 3174 2407
rect 3185 2402 3254 2407
rect 1617 2397 1622 2402
rect 1113 2392 1414 2397
rect 1425 2392 1622 2397
rect 1633 2392 1894 2397
rect 1929 2392 2142 2397
rect 2153 2392 2182 2397
rect 2177 2387 2182 2392
rect 2241 2392 2438 2397
rect 2449 2392 2630 2397
rect 2689 2392 2766 2397
rect 2785 2392 2926 2397
rect 2953 2392 3014 2397
rect 3049 2392 3126 2397
rect 3169 2392 3174 2402
rect 3185 2392 3262 2397
rect 2241 2387 2246 2392
rect 385 2382 510 2387
rect 665 2382 1030 2387
rect 1089 2382 1158 2387
rect 1201 2382 1446 2387
rect 1577 2382 1718 2387
rect 1737 2382 1974 2387
rect 2177 2382 2246 2387
rect 2265 2382 2430 2387
rect 2465 2382 2590 2387
rect 2617 2382 3086 2387
rect 3209 2382 3254 2387
rect 1577 2377 1582 2382
rect 761 2372 790 2377
rect 1121 2372 1430 2377
rect 1473 2372 1582 2377
rect 1713 2377 1718 2382
rect 2465 2377 2470 2382
rect 1713 2372 1870 2377
rect 2273 2372 2470 2377
rect 2481 2372 2902 2377
rect 2985 2372 3022 2377
rect 785 2367 1006 2372
rect 1121 2367 1126 2372
rect 1473 2367 1478 2372
rect 1001 2362 1126 2367
rect 1153 2362 1478 2367
rect 1601 2362 1870 2367
rect 2369 2362 2494 2367
rect 2545 2362 2814 2367
rect 2873 2362 2974 2367
rect 809 2352 918 2357
rect 1145 2352 1206 2357
rect 1257 2352 2206 2357
rect 2281 2352 2534 2357
rect 2609 2352 2646 2357
rect 2681 2352 2742 2357
rect 2809 2352 2870 2357
rect 2929 2352 2966 2357
rect 2609 2347 2614 2352
rect 857 2342 982 2347
rect 1177 2342 1774 2347
rect 1785 2342 1934 2347
rect 2321 2342 2374 2347
rect 2465 2342 2614 2347
rect 2641 2342 2734 2347
rect 2769 2342 3150 2347
rect 3329 2342 3358 2347
rect 633 2332 726 2337
rect 1089 2332 1126 2337
rect 1185 2332 1438 2337
rect 1561 2332 1678 2337
rect 1833 2332 1926 2337
rect 2217 2332 2302 2337
rect 2409 2332 2574 2337
rect 2793 2332 2854 2337
rect 2865 2332 2942 2337
rect 3249 2332 3366 2337
rect 865 2327 1022 2332
rect 2217 2327 2222 2332
rect 89 2322 870 2327
rect 1017 2322 1246 2327
rect 1297 2322 1646 2327
rect 1713 2322 1814 2327
rect 1713 2317 1718 2322
rect 601 2312 718 2317
rect 857 2312 1718 2317
rect 1809 2317 1814 2322
rect 1977 2322 2174 2327
rect 2193 2322 2222 2327
rect 2297 2327 2302 2332
rect 2593 2327 2774 2332
rect 2297 2322 2598 2327
rect 2769 2322 3030 2327
rect 3065 2322 3230 2327
rect 1977 2317 1982 2322
rect 1809 2312 1982 2317
rect 2169 2317 2174 2322
rect 3065 2317 3070 2322
rect 2169 2312 2334 2317
rect 2393 2312 2470 2317
rect 2513 2312 3070 2317
rect 3225 2317 3230 2322
rect 3225 2312 3254 2317
rect 3297 2312 3382 2317
rect 897 2302 1190 2307
rect 1201 2302 1318 2307
rect 1401 2302 1478 2307
rect 1729 2302 1878 2307
rect 2017 2302 2102 2307
rect 2121 2302 2278 2307
rect 2441 2302 2582 2307
rect 2817 2302 2870 2307
rect 2921 2302 2982 2307
rect 3065 2302 3134 2307
rect 3185 2302 3270 2307
rect 1537 2297 1710 2302
rect 2017 2297 2022 2302
rect 537 2292 558 2297
rect 617 2292 782 2297
rect 1041 2292 1334 2297
rect 1513 2292 1542 2297
rect 1705 2292 1790 2297
rect 1993 2292 2022 2297
rect 2097 2297 2102 2302
rect 2273 2297 2446 2302
rect 2705 2297 2822 2302
rect 2977 2297 3070 2302
rect 2097 2292 2142 2297
rect 2225 2292 2254 2297
rect 2465 2292 2550 2297
rect 2609 2292 2710 2297
rect 2841 2292 2958 2297
rect 3305 2292 3350 2297
rect 617 2287 622 2292
rect 433 2282 526 2287
rect 593 2282 622 2287
rect 777 2287 782 2292
rect 905 2287 1022 2292
rect 1329 2287 1494 2292
rect 1809 2287 1942 2292
rect 2137 2287 2230 2292
rect 2465 2287 2470 2292
rect 3097 2287 3286 2292
rect 777 2282 806 2287
rect 881 2282 910 2287
rect 1017 2282 1198 2287
rect 1217 2282 1318 2287
rect 1489 2282 1814 2287
rect 1937 2282 2118 2287
rect 2289 2282 2470 2287
rect 2673 2282 2830 2287
rect 2969 2282 3102 2287
rect 3281 2282 3374 2287
rect 521 2277 598 2282
rect 1217 2277 1222 2282
rect 2825 2277 2974 2282
rect 633 2272 1222 2277
rect 1265 2272 1670 2277
rect 1713 2272 1990 2277
rect 2225 2272 2318 2277
rect 2345 2272 2566 2277
rect 2585 2272 2694 2277
rect 3113 2272 3406 2277
rect 1665 2267 1670 2272
rect 2025 2267 2198 2272
rect 481 2262 614 2267
rect 785 2262 1646 2267
rect 1665 2262 2030 2267
rect 2193 2262 2286 2267
rect 2337 2262 2422 2267
rect 481 2257 486 2262
rect 609 2257 766 2262
rect 2561 2257 2566 2272
rect 2657 2262 2686 2267
rect 2825 2262 2950 2267
rect 3025 2262 3094 2267
rect 3241 2262 3342 2267
rect 2657 2257 2662 2262
rect 3025 2257 3030 2262
rect 3089 2257 3222 2262
rect 457 2252 486 2257
rect 761 2252 1230 2257
rect 1241 2252 1566 2257
rect 1785 2252 2038 2257
rect 2089 2252 2158 2257
rect 2177 2252 2478 2257
rect 2561 2252 2662 2257
rect 2737 2252 2894 2257
rect 3001 2252 3030 2257
rect 3217 2252 3270 2257
rect 1561 2247 1790 2252
rect 393 2242 766 2247
rect 801 2242 1006 2247
rect 1025 2242 1166 2247
rect 1257 2242 1334 2247
rect 1353 2242 1542 2247
rect 1809 2242 1918 2247
rect 2017 2242 2086 2247
rect 2129 2242 2454 2247
rect 2785 2242 2814 2247
rect 2849 2242 3286 2247
rect 1025 2237 1030 2242
rect 1913 2237 2022 2242
rect 2081 2237 2086 2242
rect 73 2232 262 2237
rect 513 2232 558 2237
rect 641 2232 1030 2237
rect 1057 2232 1710 2237
rect 1777 2232 1846 2237
rect 1857 2232 1894 2237
rect 2081 2232 2150 2237
rect 2233 2232 2302 2237
rect 2409 2232 2646 2237
rect 2665 2232 2846 2237
rect 3185 2232 3294 2237
rect 289 2222 846 2227
rect 873 2222 918 2227
rect 929 2222 1590 2227
rect 1601 2222 1718 2227
rect 1729 2222 1958 2227
rect 2265 2222 2398 2227
rect 913 2217 918 2222
rect 2641 2217 2646 2232
rect 2697 2222 2838 2227
rect 3025 2222 3166 2227
rect 3177 2222 3262 2227
rect 3329 2222 3366 2227
rect 241 2212 406 2217
rect 529 2212 902 2217
rect 913 2212 942 2217
rect 1057 2212 1246 2217
rect 1433 2212 1542 2217
rect 1569 2212 1654 2217
rect 1665 2212 2070 2217
rect 2081 2212 2174 2217
rect 2241 2212 2542 2217
rect 2641 2212 2662 2217
rect 2681 2212 2742 2217
rect 2769 2212 2814 2217
rect 2873 2212 2982 2217
rect 3065 2212 3246 2217
rect 3321 2212 3358 2217
rect 937 2207 1062 2212
rect 1265 2207 1366 2212
rect 2081 2207 2086 2212
rect 121 2202 222 2207
rect 241 2197 246 2207
rect 329 2202 590 2207
rect 785 2202 814 2207
rect 849 2202 886 2207
rect 1081 2202 1270 2207
rect 1361 2202 1766 2207
rect 1793 2202 2086 2207
rect 2097 2202 2142 2207
rect 2209 2202 2646 2207
rect 609 2197 766 2202
rect 2209 2197 2214 2202
rect 2657 2197 2662 2212
rect 2977 2207 2982 2212
rect 2713 2202 2790 2207
rect 2785 2197 2790 2202
rect 2977 2202 3006 2207
rect 185 2192 358 2197
rect 369 2192 614 2197
rect 761 2192 894 2197
rect 1001 2192 1510 2197
rect 1521 2192 1638 2197
rect 1729 2192 1982 2197
rect 2073 2192 2214 2197
rect 2233 2192 2438 2197
rect 2481 2192 2518 2197
rect 2577 2192 2598 2197
rect 2657 2192 2758 2197
rect 2785 2192 2806 2197
rect 2825 2192 2910 2197
rect 2977 2192 2982 2202
rect 3001 2197 3006 2202
rect 3105 2202 3182 2207
rect 3105 2197 3110 2202
rect 3001 2192 3110 2197
rect 3129 2192 3358 2197
rect 353 2187 358 2192
rect 209 2182 342 2187
rect 353 2182 462 2187
rect 545 2182 654 2187
rect 689 2182 1038 2187
rect 1089 2182 1134 2187
rect 1161 2182 1406 2187
rect 1417 2182 1614 2187
rect 1657 2182 2126 2187
rect 2145 2182 2614 2187
rect 3289 2182 3334 2187
rect 337 2177 342 2182
rect 545 2177 550 2182
rect 337 2172 550 2177
rect 569 2172 694 2177
rect 689 2167 694 2172
rect 817 2172 1046 2177
rect 1177 2172 1254 2177
rect 1265 2172 1686 2177
rect 1697 2172 1894 2177
rect 1929 2172 1982 2177
rect 2097 2172 2134 2177
rect 2265 2172 2550 2177
rect 817 2167 822 2172
rect 1681 2167 1686 2172
rect 2609 2167 2614 2182
rect 2625 2172 2678 2177
rect 2761 2172 2822 2177
rect 3137 2172 3366 2177
rect 385 2162 670 2167
rect 689 2162 822 2167
rect 897 2162 950 2167
rect 1081 2162 1534 2167
rect 1553 2162 1606 2167
rect 1617 2162 1654 2167
rect 1681 2162 2014 2167
rect 2057 2162 2134 2167
rect 2217 2162 2374 2167
rect 2409 2162 2462 2167
rect 2481 2162 2566 2167
rect 2609 2162 2670 2167
rect 2721 2162 2774 2167
rect 2833 2162 2926 2167
rect 3193 2162 3262 2167
rect 969 2157 1046 2162
rect 1553 2157 1558 2162
rect 2481 2157 2486 2162
rect 2833 2157 2838 2162
rect 97 2152 190 2157
rect 241 2152 294 2157
rect 481 2152 550 2157
rect 561 2152 670 2157
rect 841 2152 974 2157
rect 1041 2152 1070 2157
rect 1161 2152 1494 2157
rect 1505 2152 1558 2157
rect 1593 2152 1926 2157
rect 1945 2152 2150 2157
rect 2305 2152 2366 2157
rect 2417 2152 2438 2157
rect 2449 2152 2486 2157
rect 2497 2152 2838 2157
rect 2849 2152 2894 2157
rect 2945 2152 3038 2157
rect 3073 2152 3134 2157
rect 3305 2152 3326 2157
rect 3337 2152 3398 2157
rect 1065 2147 1166 2152
rect 137 2142 478 2147
rect 521 2142 558 2147
rect 609 2142 806 2147
rect 881 2142 902 2147
rect 913 2142 1030 2147
rect 1185 2142 1238 2147
rect 1249 2142 1358 2147
rect 1425 2142 1782 2147
rect 1817 2142 1886 2147
rect 897 2137 902 2142
rect 1233 2137 1238 2142
rect 265 2132 326 2137
rect 505 2132 702 2137
rect 897 2132 950 2137
rect 993 2132 1214 2137
rect 1233 2132 1390 2137
rect 121 2122 206 2127
rect 233 2122 302 2127
rect 425 2122 486 2127
rect 505 2122 510 2132
rect 593 2122 694 2127
rect 785 2122 1206 2127
rect 1273 2122 1318 2127
rect 1425 2122 1430 2142
rect 1521 2132 1862 2137
rect 1881 2132 1886 2142
rect 1921 2137 1926 2152
rect 2305 2147 2310 2152
rect 2449 2147 2454 2152
rect 1961 2142 2262 2147
rect 2289 2142 2310 2147
rect 2377 2142 2454 2147
rect 1921 2132 1998 2137
rect 2009 2132 2062 2137
rect 2081 2132 2398 2137
rect 2409 2132 2486 2137
rect 2513 2127 2518 2152
rect 2945 2147 2950 2152
rect 2569 2142 2814 2147
rect 2825 2142 2950 2147
rect 3033 2147 3038 2152
rect 3033 2142 3062 2147
rect 3121 2142 3222 2147
rect 3313 2142 3382 2147
rect 2553 2132 2646 2137
rect 2657 2132 3046 2137
rect 3153 2132 3230 2137
rect 121 2117 126 2122
rect 97 2112 126 2117
rect 201 2117 206 2122
rect 785 2117 790 2122
rect 1353 2117 1430 2122
rect 1465 2117 1646 2122
rect 1665 2117 1670 2127
rect 1729 2122 1838 2127
rect 1849 2122 2518 2127
rect 2545 2122 2638 2127
rect 2825 2122 3142 2127
rect 2681 2117 2774 2122
rect 201 2112 390 2117
rect 489 2112 606 2117
rect 625 2112 790 2117
rect 825 2112 950 2117
rect 993 2112 1110 2117
rect 1169 2112 1358 2117
rect 1441 2112 1470 2117
rect 1641 2112 1670 2117
rect 1729 2112 2382 2117
rect 2401 2112 2518 2117
rect 2569 2112 2646 2117
rect 2657 2112 2686 2117
rect 2769 2112 2958 2117
rect 3025 2112 3110 2117
rect 3137 2107 3142 2122
rect 3313 2112 3318 2142
rect 129 2102 190 2107
rect 273 2102 334 2107
rect 361 2102 478 2107
rect 585 2102 1214 2107
rect 1369 2102 1774 2107
rect 1785 2102 1878 2107
rect 2033 2102 2758 2107
rect 2849 2102 2910 2107
rect 2937 2102 3118 2107
rect 3137 2102 3350 2107
rect 1209 2097 1374 2102
rect 1897 2097 1982 2102
rect 2753 2097 2854 2102
rect 425 2092 566 2097
rect 593 2092 838 2097
rect 905 2092 1174 2097
rect 1393 2092 1454 2097
rect 1529 2092 1606 2097
rect 1617 2092 1902 2097
rect 1977 2092 2094 2097
rect 2121 2092 2214 2097
rect 2241 2092 2302 2097
rect 2353 2092 2486 2097
rect 2521 2092 2598 2097
rect 2617 2092 2710 2097
rect 2873 2092 2902 2097
rect 2241 2087 2246 2092
rect 2897 2087 2902 2092
rect 3097 2092 3158 2097
rect 3097 2087 3102 2092
rect 249 2082 398 2087
rect 457 2082 926 2087
rect 937 2082 1046 2087
rect 1193 2082 1342 2087
rect 1361 2082 1542 2087
rect 1633 2082 1966 2087
rect 2065 2082 2118 2087
rect 2145 2082 2246 2087
rect 2257 2082 2542 2087
rect 2561 2082 2702 2087
rect 2745 2082 2814 2087
rect 2897 2082 3102 2087
rect 249 2077 254 2082
rect 225 2072 254 2077
rect 393 2077 398 2082
rect 1041 2077 1046 2082
rect 1065 2077 1198 2082
rect 1337 2077 1342 2082
rect 393 2072 422 2077
rect 433 2072 526 2077
rect 657 2072 1022 2077
rect 1041 2072 1070 2077
rect 1337 2072 1646 2077
rect 1697 2072 1766 2077
rect 1857 2072 1958 2077
rect 1969 2072 1990 2077
rect 2041 2072 2102 2077
rect 2177 2072 2438 2077
rect 2473 2072 2582 2077
rect 2593 2072 2830 2077
rect 545 2067 662 2072
rect 1217 2067 1318 2072
rect 153 2062 550 2067
rect 673 2062 846 2067
rect 865 2062 886 2067
rect 897 2062 1222 2067
rect 1313 2062 1838 2067
rect 1905 2062 2038 2067
rect 2265 2062 2374 2067
rect 2161 2057 2246 2062
rect 2433 2057 2438 2072
rect 2449 2062 2774 2067
rect 2785 2062 2982 2067
rect 337 2052 478 2057
rect 505 2052 1134 2057
rect 1177 2052 1222 2057
rect 1265 2052 2166 2057
rect 2241 2052 2406 2057
rect 2433 2052 2598 2057
rect 2609 2052 2654 2057
rect 2665 2052 2894 2057
rect 241 2047 318 2052
rect 2913 2047 3006 2052
rect 161 2042 246 2047
rect 313 2042 358 2047
rect 401 2042 430 2047
rect 537 2042 566 2047
rect 649 2042 902 2047
rect 953 2042 1006 2047
rect 1025 2042 1446 2047
rect 1553 2042 1654 2047
rect 1681 2042 1790 2047
rect 1921 2042 1990 2047
rect 2177 2042 2478 2047
rect 2505 2042 2726 2047
rect 2801 2042 2918 2047
rect 3001 2042 3030 2047
rect 3161 2042 3262 2047
rect 425 2037 542 2042
rect 2801 2037 2806 2042
rect 257 2032 382 2037
rect 561 2032 630 2037
rect 665 2032 718 2037
rect 737 2032 1230 2037
rect 1289 2032 1366 2037
rect 1441 2032 1478 2037
rect 1497 2032 1630 2037
rect 1641 2032 1862 2037
rect 1873 2032 2038 2037
rect 2073 2032 2142 2037
rect 2233 2032 2462 2037
rect 2473 2032 2806 2037
rect 2817 2032 2990 2037
rect 3081 2032 3150 2037
rect 561 2027 566 2032
rect 2033 2027 2038 2032
rect 3145 2027 3150 2032
rect 3273 2032 3382 2037
rect 3273 2027 3278 2032
rect 169 2022 254 2027
rect 345 2022 438 2027
rect 481 2022 566 2027
rect 585 2022 918 2027
rect 945 2022 1558 2027
rect 1665 2022 2022 2027
rect 2033 2022 2182 2027
rect 2297 2022 2326 2027
rect 2361 2022 2422 2027
rect 2441 2022 2710 2027
rect 2721 2022 2942 2027
rect 2953 2022 3102 2027
rect 3145 2022 3278 2027
rect 2017 2017 2022 2022
rect 393 2012 822 2017
rect 833 2012 1438 2017
rect 1593 2012 2006 2017
rect 2017 2012 2278 2017
rect 2289 2012 2582 2017
rect 2905 2012 3014 2017
rect 2601 2007 2886 2012
rect 177 2002 310 2007
rect 329 2002 638 2007
rect 681 2002 1030 2007
rect 1257 2002 1518 2007
rect 1553 2002 1574 2007
rect 1609 2002 1638 2007
rect 1761 2002 1798 2007
rect 1873 2002 1942 2007
rect 1969 2002 2606 2007
rect 2881 2002 3110 2007
rect 305 1997 310 2002
rect 1049 1997 1230 2002
rect 65 1992 286 1997
rect 305 1992 982 1997
rect 1001 1992 1054 1997
rect 1225 1992 1254 1997
rect 1273 1992 1334 1997
rect 1401 1992 2390 1997
rect 2409 1992 2470 1997
rect 2545 1992 3150 1997
rect 3217 1992 3318 1997
rect 977 1987 982 1992
rect 81 1982 382 1987
rect 457 1982 694 1987
rect 713 1982 774 1987
rect 785 1982 806 1987
rect 865 1982 894 1987
rect 913 1982 950 1987
rect 977 1982 1502 1987
rect 1545 1982 1574 1987
rect 1593 1982 1862 1987
rect 1961 1982 2230 1987
rect 2241 1982 2846 1987
rect 2857 1982 2942 1987
rect 2969 1982 3046 1987
rect 3073 1982 3238 1987
rect 3265 1982 3310 1987
rect 769 1977 774 1982
rect 1569 1977 1574 1982
rect 153 1972 230 1977
rect 385 1972 574 1977
rect 729 1972 758 1977
rect 769 1972 950 1977
rect 969 1972 1246 1977
rect 1257 1972 1558 1977
rect 1569 1972 1654 1977
rect 1689 1972 1782 1977
rect 1793 1972 1838 1977
rect 249 1967 366 1972
rect 569 1967 734 1972
rect 1553 1967 1558 1972
rect 1857 1967 1862 1982
rect 3041 1977 3046 1982
rect 1897 1972 1958 1977
rect 2017 1972 2062 1977
rect 2073 1972 2110 1977
rect 2121 1972 2198 1977
rect 2265 1972 2318 1977
rect 2353 1972 2654 1977
rect 2681 1972 2806 1977
rect 2817 1972 3014 1977
rect 3041 1972 3150 1977
rect 2801 1967 2806 1972
rect 3169 1967 3262 1972
rect 193 1962 254 1967
rect 361 1962 414 1967
rect 481 1962 550 1967
rect 769 1962 1302 1967
rect 1329 1962 1358 1967
rect 1409 1962 1486 1967
rect 1553 1962 1846 1967
rect 1857 1962 1998 1967
rect 2009 1962 2254 1967
rect 2313 1962 2342 1967
rect 2433 1962 2478 1967
rect 2505 1962 2614 1967
rect 2625 1962 2766 1967
rect 2801 1962 2894 1967
rect 2905 1962 3174 1967
rect 3257 1962 3286 1967
rect 2433 1957 2438 1962
rect 2609 1957 2614 1962
rect 113 1952 166 1957
rect 241 1952 270 1957
rect 313 1952 470 1957
rect 513 1952 566 1957
rect 593 1952 646 1957
rect 657 1952 686 1957
rect 705 1952 990 1957
rect 1001 1952 1054 1957
rect 1153 1952 1222 1957
rect 1233 1952 1390 1957
rect 1473 1952 1686 1957
rect 1713 1952 1782 1957
rect 1817 1952 1886 1957
rect 1953 1952 2046 1957
rect 2105 1952 2166 1957
rect 2177 1952 2198 1957
rect 2225 1952 2438 1957
rect 2457 1952 2550 1957
rect 2609 1952 2734 1957
rect 2937 1952 3030 1957
rect 1217 1947 1222 1952
rect 1385 1947 1478 1952
rect 1777 1947 1782 1952
rect 2177 1947 2182 1952
rect 3161 1947 3166 1957
rect 3185 1952 3254 1957
rect 65 1942 110 1947
rect 161 1942 190 1947
rect 297 1942 662 1947
rect 713 1942 814 1947
rect 841 1942 1198 1947
rect 1217 1942 1270 1947
rect 1289 1942 1366 1947
rect 1497 1942 1702 1947
rect 1745 1942 1766 1947
rect 1777 1942 2302 1947
rect 2337 1942 2470 1947
rect 2529 1942 2630 1947
rect 2641 1942 2694 1947
rect 65 1917 70 1942
rect 89 1932 134 1937
rect 161 1927 166 1942
rect 657 1937 662 1942
rect 1745 1937 1750 1942
rect 2465 1937 2470 1942
rect 113 1922 166 1927
rect 177 1927 182 1937
rect 193 1932 230 1937
rect 265 1932 374 1937
rect 441 1932 462 1937
rect 489 1932 606 1937
rect 657 1932 974 1937
rect 1065 1932 1510 1937
rect 1569 1932 1726 1937
rect 1745 1932 1760 1937
rect 1769 1932 1838 1937
rect 1857 1932 1918 1937
rect 1937 1932 1990 1937
rect 2081 1932 2166 1937
rect 2209 1932 2326 1937
rect 2361 1932 2454 1937
rect 2465 1932 2686 1937
rect 177 1922 238 1927
rect 257 1922 350 1927
rect 369 1922 374 1932
rect 1755 1927 1760 1932
rect 401 1922 446 1927
rect 473 1922 518 1927
rect 529 1922 862 1927
rect 905 1922 1078 1927
rect 1161 1922 1518 1927
rect 1537 1922 1598 1927
rect 1697 1922 1750 1927
rect 1755 1922 1782 1927
rect 417 1917 422 1922
rect 1073 1917 1166 1922
rect 1537 1917 1542 1922
rect 1793 1917 1798 1927
rect 65 1912 110 1917
rect 217 1912 286 1917
rect 417 1912 502 1917
rect 513 1912 734 1917
rect 745 1912 814 1917
rect 993 1912 1014 1917
rect 1185 1912 1254 1917
rect 1313 1912 1542 1917
rect 1601 1912 1798 1917
rect 1809 1912 1846 1917
rect 1857 1912 1862 1932
rect 2161 1927 2166 1932
rect 2705 1927 2710 1947
rect 2745 1942 2774 1947
rect 2833 1942 2926 1947
rect 2993 1942 3142 1947
rect 3153 1942 3166 1947
rect 3177 1942 3262 1947
rect 2921 1937 2998 1942
rect 3153 1937 3158 1942
rect 2785 1927 2790 1937
rect 2825 1932 2870 1937
rect 2865 1927 2870 1932
rect 2081 1922 2102 1927
rect 2111 1922 2142 1927
rect 2161 1922 2190 1927
rect 2081 1917 2086 1922
rect 1873 1912 1910 1917
rect 1985 1912 2086 1917
rect 161 1902 294 1907
rect 313 1902 350 1907
rect 377 1902 470 1907
rect 513 1902 518 1912
rect 849 1907 974 1912
rect 1313 1907 1318 1912
rect 2111 1907 2116 1922
rect 2185 1917 2190 1922
rect 2249 1922 2326 1927
rect 2433 1922 2534 1927
rect 2561 1922 2646 1927
rect 2665 1922 2710 1927
rect 2753 1922 2790 1927
rect 2841 1922 2870 1927
rect 2249 1917 2254 1922
rect 2121 1912 2166 1917
rect 2185 1912 2254 1917
rect 609 1902 638 1907
rect 657 1902 686 1907
rect 753 1902 854 1907
rect 969 1902 1318 1907
rect 1337 1902 1406 1907
rect 1457 1902 1502 1907
rect 1633 1902 1918 1907
rect 2017 1902 2062 1907
rect 2081 1902 2116 1907
rect 1521 1897 1614 1902
rect 169 1892 190 1897
rect 233 1892 406 1897
rect 481 1892 574 1897
rect 593 1892 654 1897
rect 673 1892 782 1897
rect 865 1892 1078 1897
rect 1137 1892 1526 1897
rect 1609 1892 1934 1897
rect 2009 1892 2110 1897
rect 2121 1892 2150 1897
rect 2161 1892 2262 1897
rect 2161 1887 2166 1892
rect 2321 1887 2326 1922
rect 2369 1912 2854 1917
rect 2881 1912 2886 1937
rect 3017 1932 3158 1937
rect 2937 1922 3062 1927
rect 3177 1922 3222 1927
rect 2929 1912 2990 1917
rect 3097 1912 3142 1917
rect 3153 1912 3190 1917
rect 3241 1912 3318 1917
rect 3241 1907 3246 1912
rect 2401 1902 2870 1907
rect 2889 1902 2958 1907
rect 3129 1902 3246 1907
rect 3313 1907 3318 1912
rect 3313 1902 3358 1907
rect 2369 1892 2974 1897
rect 3193 1892 3302 1897
rect 361 1882 686 1887
rect 913 1882 1094 1887
rect 1337 1882 1382 1887
rect 1441 1882 1694 1887
rect 1801 1882 2166 1887
rect 2185 1882 2286 1887
rect 2321 1882 2518 1887
rect 2529 1882 2590 1887
rect 2617 1882 2694 1887
rect 2705 1882 2822 1887
rect 2833 1882 3038 1887
rect 3153 1882 3254 1887
rect 1129 1877 1318 1882
rect 3153 1877 3158 1882
rect 81 1872 422 1877
rect 545 1872 630 1877
rect 673 1872 742 1877
rect 1105 1872 1134 1877
rect 1313 1872 1398 1877
rect 1417 1872 1462 1877
rect 1529 1872 1566 1877
rect 1641 1872 1702 1877
rect 1753 1872 1870 1877
rect 2097 1872 2174 1877
rect 2377 1872 2462 1877
rect 2481 1872 2542 1877
rect 2593 1872 2622 1877
rect 2697 1872 2790 1877
rect 2801 1872 2838 1877
rect 2849 1872 3022 1877
rect 3057 1872 3158 1877
rect 993 1867 1086 1872
rect 1393 1867 1398 1872
rect 1889 1867 2078 1872
rect 2785 1867 2790 1872
rect 3057 1867 3062 1872
rect 257 1862 582 1867
rect 761 1862 894 1867
rect 969 1862 998 1867
rect 1081 1862 1366 1867
rect 1393 1862 1438 1867
rect 1497 1862 1894 1867
rect 2073 1862 2230 1867
rect 2321 1862 2350 1867
rect 2441 1862 2710 1867
rect 2785 1862 3062 1867
rect 3201 1862 3238 1867
rect 113 1852 150 1857
rect 145 1842 246 1847
rect 129 1807 134 1837
rect 113 1802 134 1807
rect 241 1807 246 1817
rect 257 1812 262 1862
rect 601 1857 766 1862
rect 889 1857 894 1862
rect 377 1852 606 1857
rect 889 1852 1190 1857
rect 1345 1852 2470 1857
rect 2537 1852 2662 1857
rect 2729 1852 3062 1857
rect 3081 1852 3230 1857
rect 289 1842 342 1847
rect 385 1842 518 1847
rect 577 1842 630 1847
rect 665 1842 702 1847
rect 1025 1842 1902 1847
rect 1937 1842 2206 1847
rect 2241 1842 2278 1847
rect 2289 1842 2406 1847
rect 2417 1842 2702 1847
rect 2777 1842 2854 1847
rect 2889 1842 3006 1847
rect 3137 1842 3254 1847
rect 721 1837 790 1842
rect 833 1837 950 1842
rect 3025 1837 3142 1842
rect 329 1832 726 1837
rect 785 1832 838 1837
rect 945 1832 1014 1837
rect 1009 1827 1014 1832
rect 1097 1832 1238 1837
rect 1497 1832 1990 1837
rect 2073 1832 2350 1837
rect 2393 1832 3030 1837
rect 3153 1832 3318 1837
rect 1097 1827 1102 1832
rect 1233 1827 1478 1832
rect 1985 1827 2078 1832
rect 3153 1827 3158 1832
rect 377 1822 438 1827
rect 489 1822 550 1827
rect 665 1822 774 1827
rect 849 1822 934 1827
rect 1009 1822 1102 1827
rect 1161 1822 1182 1827
rect 1473 1822 1510 1827
rect 1537 1822 1566 1827
rect 1577 1822 1966 1827
rect 2097 1822 2142 1827
rect 2153 1822 2246 1827
rect 2257 1822 2294 1827
rect 2361 1822 2446 1827
rect 2457 1822 2558 1827
rect 2577 1822 2774 1827
rect 2785 1822 2814 1827
rect 2913 1822 3086 1827
rect 3129 1822 3158 1827
rect 3177 1822 3310 1827
rect 273 1807 278 1817
rect 337 1812 366 1817
rect 409 1812 446 1817
rect 465 1812 518 1817
rect 745 1812 870 1817
rect 1161 1812 1374 1817
rect 1433 1812 1614 1817
rect 1697 1812 1838 1817
rect 1913 1812 2990 1817
rect 3209 1812 3326 1817
rect 241 1802 278 1807
rect 401 1802 502 1807
rect 401 1797 406 1802
rect 513 1797 518 1812
rect 537 1802 742 1807
rect 769 1802 830 1807
rect 849 1802 902 1807
rect 913 1802 1030 1807
rect 1161 1802 1166 1812
rect 3009 1807 3158 1812
rect 1209 1802 1438 1807
rect 1553 1802 1990 1807
rect 2065 1802 2278 1807
rect 2345 1802 2590 1807
rect 2633 1802 2910 1807
rect 2953 1802 3014 1807
rect 3153 1802 3198 1807
rect 3265 1802 3310 1807
rect 849 1797 854 1802
rect 3193 1797 3270 1802
rect 169 1792 350 1797
rect 385 1792 430 1797
rect 513 1792 542 1797
rect 553 1792 590 1797
rect 825 1792 854 1797
rect 1049 1792 1142 1797
rect 1225 1792 1502 1797
rect 1521 1792 1582 1797
rect 1697 1792 2302 1797
rect 2329 1792 2390 1797
rect 2449 1792 3142 1797
rect 3289 1792 3334 1797
rect 1049 1787 1054 1792
rect 105 1782 190 1787
rect 249 1782 342 1787
rect 401 1777 406 1787
rect 417 1782 550 1787
rect 609 1782 806 1787
rect 929 1782 1054 1787
rect 1137 1787 1142 1792
rect 1137 1782 1726 1787
rect 1745 1782 1974 1787
rect 1985 1782 2038 1787
rect 2057 1782 2214 1787
rect 2257 1782 2502 1787
rect 2553 1782 2726 1787
rect 2737 1782 2942 1787
rect 2993 1782 3134 1787
rect 3201 1782 3350 1787
rect 417 1777 422 1782
rect 609 1777 614 1782
rect 329 1772 406 1777
rect 409 1772 422 1777
rect 497 1772 614 1777
rect 801 1777 806 1782
rect 2721 1777 2726 1782
rect 801 1772 878 1777
rect 1049 1772 1470 1777
rect 1537 1772 1622 1777
rect 1665 1772 2126 1777
rect 2177 1772 2214 1777
rect 2225 1772 2470 1777
rect 2481 1772 2502 1777
rect 2513 1772 2670 1777
rect 2721 1772 2918 1777
rect 2969 1772 2998 1777
rect 3073 1772 3110 1777
rect 3161 1772 3398 1777
rect 409 1767 414 1772
rect 2209 1767 2214 1772
rect 2465 1767 2470 1772
rect 2497 1767 2502 1772
rect 2913 1767 2918 1772
rect 233 1762 414 1767
rect 497 1762 598 1767
rect 609 1762 886 1767
rect 1009 1762 1302 1767
rect 1337 1762 1646 1767
rect 1737 1762 1822 1767
rect 1833 1762 1878 1767
rect 1937 1762 2142 1767
rect 2209 1762 2262 1767
rect 2321 1762 2454 1767
rect 2465 1762 2486 1767
rect 2497 1762 2686 1767
rect 2729 1762 2814 1767
rect 2913 1762 3030 1767
rect 3049 1762 3086 1767
rect 3105 1762 3190 1767
rect 3209 1762 3238 1767
rect 3185 1757 3190 1762
rect 3297 1757 3302 1767
rect 353 1752 470 1757
rect 601 1752 630 1757
rect 737 1752 998 1757
rect 1129 1752 1662 1757
rect 1953 1752 2118 1757
rect 2145 1752 2166 1757
rect 2185 1752 2478 1757
rect 2505 1752 2574 1757
rect 2625 1752 2814 1757
rect 2937 1752 2958 1757
rect 2969 1752 3102 1757
rect 3185 1752 3302 1757
rect 625 1747 742 1752
rect 993 1747 1134 1752
rect 65 1742 86 1747
rect 113 1742 182 1747
rect 233 1742 254 1747
rect 449 1742 534 1747
rect 553 1742 590 1747
rect 761 1742 790 1747
rect 81 1707 86 1742
rect 785 1737 790 1742
rect 865 1742 894 1747
rect 1369 1742 1590 1747
rect 1625 1742 1662 1747
rect 1681 1742 1774 1747
rect 1793 1742 1814 1747
rect 1929 1742 2014 1747
rect 2041 1742 2174 1747
rect 2297 1742 2358 1747
rect 2417 1742 2446 1747
rect 2457 1742 2662 1747
rect 2689 1742 2726 1747
rect 2737 1742 2806 1747
rect 2873 1742 2910 1747
rect 2953 1742 3054 1747
rect 3201 1742 3246 1747
rect 865 1737 870 1742
rect 1793 1737 1798 1742
rect 97 1712 102 1737
rect 129 1732 158 1737
rect 201 1732 230 1737
rect 265 1732 310 1737
rect 337 1732 550 1737
rect 569 1732 654 1737
rect 697 1732 742 1737
rect 785 1732 870 1737
rect 1065 1732 1182 1737
rect 1273 1732 1398 1737
rect 1497 1732 1798 1737
rect 1817 1732 2710 1737
rect 81 1702 118 1707
rect 129 1697 134 1732
rect 225 1727 230 1732
rect 185 1722 230 1727
rect 329 1722 430 1727
rect 529 1722 582 1727
rect 633 1722 702 1727
rect 1137 1722 1238 1727
rect 1321 1722 1574 1727
rect 1633 1722 2054 1727
rect 2065 1722 2158 1727
rect 2241 1722 2366 1727
rect 2409 1722 2470 1727
rect 2585 1722 2662 1727
rect 529 1717 534 1722
rect 1233 1717 1238 1722
rect 2465 1717 2470 1722
rect 193 1712 246 1717
rect 281 1712 342 1717
rect 417 1712 462 1717
rect 529 1712 558 1717
rect 577 1712 598 1717
rect 641 1712 846 1717
rect 953 1712 974 1717
rect 1137 1712 1222 1717
rect 1233 1712 1366 1717
rect 1377 1712 1398 1717
rect 1425 1712 1710 1717
rect 1825 1712 2374 1717
rect 2465 1712 2550 1717
rect 2569 1712 2622 1717
rect 2641 1712 2694 1717
rect 1705 1707 1830 1712
rect 2545 1707 2550 1712
rect 2705 1707 2710 1732
rect 2721 1717 2726 1742
rect 3073 1737 3182 1742
rect 2737 1732 2774 1737
rect 2793 1732 2830 1737
rect 2841 1732 3078 1737
rect 3177 1732 3310 1737
rect 2737 1722 2742 1732
rect 2769 1717 2774 1732
rect 2825 1722 2830 1732
rect 2849 1722 3278 1727
rect 3345 1722 3398 1727
rect 2721 1712 2758 1717
rect 2769 1712 2822 1717
rect 2833 1712 2886 1717
rect 2953 1712 3046 1717
rect 3057 1712 3198 1717
rect 3041 1707 3046 1712
rect 153 1702 238 1707
rect 281 1702 310 1707
rect 321 1702 342 1707
rect 521 1702 1022 1707
rect 1041 1702 1310 1707
rect 1369 1702 1518 1707
rect 1529 1702 1686 1707
rect 2001 1702 2062 1707
rect 2137 1702 2446 1707
rect 2545 1702 2662 1707
rect 2705 1702 2862 1707
rect 2889 1702 3030 1707
rect 3041 1702 3062 1707
rect 3097 1702 3374 1707
rect 1041 1697 1046 1702
rect 1849 1697 1926 1702
rect 65 1692 134 1697
rect 161 1692 206 1697
rect 249 1692 278 1697
rect 353 1692 1046 1697
rect 1129 1692 1214 1697
rect 1489 1692 1854 1697
rect 1921 1692 2550 1697
rect 2577 1692 2614 1697
rect 2625 1692 2734 1697
rect 2825 1692 3158 1697
rect 3201 1692 3246 1697
rect 65 1677 70 1692
rect 273 1687 358 1692
rect 1289 1687 1470 1692
rect 2545 1687 2550 1692
rect 81 1682 126 1687
rect 145 1682 166 1687
rect 537 1682 1150 1687
rect 1225 1682 1294 1687
rect 1465 1682 1510 1687
rect 1593 1682 1686 1687
rect 1865 1682 1910 1687
rect 2025 1682 2110 1687
rect 2209 1682 2302 1687
rect 2449 1682 2534 1687
rect 2545 1682 3070 1687
rect 3145 1682 3174 1687
rect 3233 1682 3294 1687
rect 417 1677 502 1682
rect 1145 1677 1230 1682
rect 2321 1677 2406 1682
rect 65 1672 158 1677
rect 305 1672 422 1677
rect 497 1672 734 1677
rect 889 1672 1126 1677
rect 1305 1672 1430 1677
rect 1441 1672 1878 1677
rect 1889 1672 2326 1677
rect 2401 1672 2438 1677
rect 2505 1672 3254 1677
rect 729 1667 894 1672
rect 1425 1667 1430 1672
rect 1873 1667 1878 1672
rect 2433 1667 2510 1672
rect 105 1662 294 1667
rect 433 1662 486 1667
rect 569 1662 606 1667
rect 625 1662 670 1667
rect 681 1662 710 1667
rect 913 1662 966 1667
rect 1129 1662 1174 1667
rect 1217 1662 1414 1667
rect 1425 1662 1502 1667
rect 1545 1662 1710 1667
rect 1873 1662 2102 1667
rect 2113 1662 2390 1667
rect 2529 1662 2598 1667
rect 2649 1662 3014 1667
rect 3025 1662 3342 1667
rect 289 1657 438 1662
rect 985 1657 1110 1662
rect 3025 1657 3030 1662
rect 457 1652 990 1657
rect 1105 1652 1206 1657
rect 1321 1652 1742 1657
rect 1857 1652 1902 1657
rect 2065 1652 2174 1657
rect 2193 1652 2254 1657
rect 2337 1652 3030 1657
rect 3057 1652 3118 1657
rect 3209 1652 3238 1657
rect 1201 1647 1326 1652
rect 2065 1647 2070 1652
rect 3113 1647 3214 1652
rect 289 1642 382 1647
rect 497 1642 1078 1647
rect 1089 1642 1182 1647
rect 1345 1642 2070 1647
rect 2089 1642 2198 1647
rect 2281 1642 2358 1647
rect 2473 1642 3094 1647
rect 497 1637 502 1642
rect 1073 1637 1078 1642
rect 105 1632 150 1637
rect 241 1632 502 1637
rect 521 1632 614 1637
rect 633 1632 1054 1637
rect 1073 1632 1286 1637
rect 1457 1632 1558 1637
rect 1601 1632 1622 1637
rect 1633 1632 1678 1637
rect 1777 1632 1902 1637
rect 2009 1632 2158 1637
rect 2241 1632 2310 1637
rect 2393 1632 3118 1637
rect 3129 1632 3262 1637
rect 3305 1632 3398 1637
rect 97 1622 118 1627
rect 177 1622 230 1627
rect 361 1622 390 1627
rect 97 1607 102 1622
rect 177 1617 182 1622
rect 249 1617 326 1622
rect 113 1612 182 1617
rect 193 1612 254 1617
rect 321 1612 518 1617
rect 97 1602 118 1607
rect 209 1602 310 1607
rect 457 1602 478 1607
rect 209 1597 214 1602
rect 73 1592 126 1597
rect 193 1592 214 1597
rect 225 1592 254 1597
rect 377 1592 502 1597
rect 513 1592 518 1612
rect 609 1597 614 1632
rect 1321 1627 1462 1632
rect 1553 1627 1558 1632
rect 681 1622 710 1627
rect 705 1617 710 1622
rect 777 1622 910 1627
rect 937 1622 1062 1627
rect 1145 1622 1246 1627
rect 1297 1622 1326 1627
rect 1481 1622 1542 1627
rect 1553 1622 1614 1627
rect 1625 1622 3182 1627
rect 777 1617 782 1622
rect 705 1612 782 1617
rect 801 1612 862 1617
rect 961 1612 1054 1617
rect 1281 1612 1414 1617
rect 1793 1612 1910 1617
rect 1937 1612 1966 1617
rect 1993 1612 2446 1617
rect 2593 1612 2718 1617
rect 2897 1612 2918 1617
rect 2969 1612 3030 1617
rect 3065 1612 3094 1617
rect 3225 1612 3262 1617
rect 3297 1612 3350 1617
rect 1073 1607 1246 1612
rect 1409 1607 1414 1612
rect 1561 1607 1630 1612
rect 1713 1607 1798 1612
rect 2145 1607 2150 1612
rect 961 1602 1078 1607
rect 1241 1602 1390 1607
rect 1409 1602 1566 1607
rect 1625 1602 1718 1607
rect 1817 1602 2006 1607
rect 2033 1602 2054 1607
rect 2065 1602 2102 1607
rect 2113 1602 2150 1607
rect 2185 1602 2358 1607
rect 2369 1602 2374 1612
rect 2441 1607 2598 1612
rect 2713 1607 2886 1612
rect 2385 1602 2422 1607
rect 2617 1602 2694 1607
rect 2881 1602 3062 1607
rect 3097 1602 3158 1607
rect 2353 1597 2358 1602
rect 609 1592 686 1597
rect 833 1592 1230 1597
rect 1345 1592 1406 1597
rect 1577 1592 1630 1597
rect 1673 1592 1726 1597
rect 1737 1592 2342 1597
rect 2353 1592 2374 1597
rect 1225 1587 1334 1592
rect 1401 1587 1582 1592
rect 2337 1587 2342 1592
rect 81 1582 126 1587
rect 193 1582 278 1587
rect 305 1582 334 1587
rect 577 1582 646 1587
rect 665 1582 694 1587
rect 913 1582 942 1587
rect 993 1582 1054 1587
rect 1073 1582 1206 1587
rect 1329 1582 1382 1587
rect 1601 1582 1622 1587
rect 1665 1582 1702 1587
rect 1737 1582 1966 1587
rect 1977 1582 2014 1587
rect 2025 1582 2102 1587
rect 2257 1582 2326 1587
rect 2337 1582 2366 1587
rect 2121 1577 2230 1582
rect 2385 1577 2390 1602
rect 2401 1592 2590 1597
rect 2633 1592 2726 1597
rect 2801 1592 3190 1597
rect 2609 1582 2670 1587
rect 2689 1582 2718 1587
rect 2865 1582 3118 1587
rect 3161 1582 3214 1587
rect 49 1572 142 1577
rect 217 1572 358 1577
rect 385 1572 502 1577
rect 561 1572 702 1577
rect 841 1572 934 1577
rect 1185 1572 1262 1577
rect 1425 1572 1494 1577
rect 1561 1572 1582 1577
rect 1633 1572 1678 1577
rect 1713 1572 2126 1577
rect 2225 1572 2390 1577
rect 2561 1572 2686 1577
rect 2785 1572 2862 1577
rect 2929 1572 3006 1577
rect 3033 1572 3142 1577
rect 3169 1572 3190 1577
rect 49 1477 54 1572
rect 929 1567 1022 1572
rect 1057 1567 1166 1572
rect 1281 1567 1366 1572
rect 1425 1567 1430 1572
rect 65 1562 134 1567
rect 177 1562 230 1567
rect 289 1562 478 1567
rect 561 1562 598 1567
rect 761 1562 910 1567
rect 1017 1562 1062 1567
rect 1161 1562 1286 1567
rect 1361 1562 1430 1567
rect 1489 1567 1494 1572
rect 1489 1562 1550 1567
rect 1665 1562 1974 1567
rect 2001 1562 2110 1567
rect 2121 1562 2214 1567
rect 2321 1562 2382 1567
rect 2457 1562 2942 1567
rect 2985 1562 3238 1567
rect 65 1487 70 1562
rect 1545 1557 1670 1562
rect 81 1552 174 1557
rect 241 1552 550 1557
rect 777 1552 894 1557
rect 953 1552 1006 1557
rect 1073 1552 1166 1557
rect 1225 1552 1350 1557
rect 1441 1552 1478 1557
rect 1689 1552 1814 1557
rect 1857 1552 1878 1557
rect 1897 1552 1926 1557
rect 1969 1552 2118 1557
rect 2169 1552 2334 1557
rect 2449 1552 2534 1557
rect 2593 1552 2734 1557
rect 2777 1552 3150 1557
rect 3273 1552 3350 1557
rect 81 1542 102 1547
rect 145 1542 278 1547
rect 305 1542 358 1547
rect 393 1542 438 1547
rect 601 1542 630 1547
rect 649 1542 742 1547
rect 857 1542 1126 1547
rect 1177 1542 1334 1547
rect 1345 1542 1414 1547
rect 81 1497 86 1542
rect 193 1532 334 1537
rect 193 1517 198 1532
rect 265 1522 318 1527
rect 137 1512 198 1517
rect 217 1512 326 1517
rect 353 1507 358 1542
rect 649 1537 654 1542
rect 737 1537 838 1542
rect 1441 1537 1446 1552
rect 1969 1547 1974 1552
rect 2529 1547 2534 1552
rect 1465 1542 1510 1547
rect 1625 1542 1862 1547
rect 1905 1542 1974 1547
rect 2033 1542 2190 1547
rect 2201 1542 2286 1547
rect 2305 1542 2334 1547
rect 2353 1542 2518 1547
rect 2529 1542 2614 1547
rect 2641 1542 2886 1547
rect 2905 1542 2958 1547
rect 3033 1542 3078 1547
rect 3089 1542 3134 1547
rect 3337 1542 3398 1547
rect 2609 1537 2614 1542
rect 369 1532 502 1537
rect 593 1532 654 1537
rect 833 1532 1014 1537
rect 1169 1532 1422 1537
rect 1441 1532 1478 1537
rect 1489 1532 1742 1537
rect 1785 1532 1806 1537
rect 1841 1532 1998 1537
rect 2017 1532 2134 1537
rect 2153 1532 2478 1537
rect 2537 1532 2590 1537
rect 2609 1532 2638 1537
rect 1033 1527 1150 1532
rect 1841 1527 1846 1532
rect 2129 1527 2134 1532
rect 2633 1527 2774 1532
rect 377 1522 422 1527
rect 441 1522 518 1527
rect 545 1522 1038 1527
rect 1145 1522 1510 1527
rect 1649 1522 1846 1527
rect 1905 1522 1942 1527
rect 2129 1522 2238 1527
rect 2265 1522 2366 1527
rect 513 1517 518 1522
rect 1649 1517 1654 1522
rect 433 1512 486 1517
rect 513 1512 1654 1517
rect 1697 1512 2030 1517
rect 2041 1512 2182 1517
rect 2201 1512 2310 1517
rect 2465 1512 2518 1517
rect 2617 1512 2726 1517
rect 2617 1507 2622 1512
rect 105 1502 134 1507
rect 185 1502 222 1507
rect 321 1502 422 1507
rect 481 1502 510 1507
rect 617 1502 766 1507
rect 817 1502 1294 1507
rect 1409 1502 1990 1507
rect 2009 1502 2062 1507
rect 2097 1502 2118 1507
rect 2137 1502 2334 1507
rect 2409 1502 2622 1507
rect 2721 1507 2726 1512
rect 2769 1507 2774 1527
rect 2817 1512 2822 1537
rect 2913 1532 3014 1537
rect 3073 1532 3126 1537
rect 3193 1532 3270 1537
rect 3281 1532 3334 1537
rect 2857 1522 2902 1527
rect 2929 1522 2990 1527
rect 3201 1522 3294 1527
rect 3345 1522 3398 1527
rect 3345 1517 3350 1522
rect 2969 1512 3038 1517
rect 3065 1512 3190 1517
rect 3209 1512 3238 1517
rect 3185 1507 3190 1512
rect 3233 1507 3238 1512
rect 3305 1512 3350 1517
rect 3305 1507 3310 1512
rect 2721 1502 2750 1507
rect 2769 1502 2998 1507
rect 3017 1502 3134 1507
rect 3185 1502 3206 1507
rect 3233 1502 3310 1507
rect 505 1497 622 1502
rect 81 1492 102 1497
rect 113 1492 246 1497
rect 641 1492 798 1497
rect 817 1487 822 1502
rect 1289 1497 1414 1502
rect 1985 1497 1990 1502
rect 2113 1497 2118 1502
rect 873 1492 902 1497
rect 953 1492 1270 1497
rect 1433 1492 1502 1497
rect 1545 1492 1614 1497
rect 1705 1492 1734 1497
rect 1729 1487 1734 1492
rect 1809 1492 1838 1497
rect 1865 1492 1918 1497
rect 1985 1492 2102 1497
rect 2113 1492 2166 1497
rect 2297 1492 2366 1497
rect 2441 1492 2526 1497
rect 2633 1492 2798 1497
rect 2953 1492 3142 1497
rect 1809 1487 1814 1492
rect 2161 1487 2302 1492
rect 65 1482 134 1487
rect 193 1482 270 1487
rect 289 1482 366 1487
rect 513 1482 734 1487
rect 761 1482 822 1487
rect 913 1482 1230 1487
rect 1313 1482 1366 1487
rect 1593 1482 1710 1487
rect 1729 1482 1814 1487
rect 2073 1482 2142 1487
rect 2553 1482 2622 1487
rect 2809 1482 2958 1487
rect 2985 1482 3006 1487
rect 3033 1482 3094 1487
rect 289 1477 294 1482
rect 49 1472 142 1477
rect 169 1472 294 1477
rect 361 1477 366 1482
rect 1385 1477 1502 1482
rect 2617 1477 2814 1482
rect 361 1472 390 1477
rect 449 1472 598 1477
rect 609 1472 638 1477
rect 961 1472 1030 1477
rect 1153 1472 1390 1477
rect 1497 1472 1598 1477
rect 1953 1472 2070 1477
rect 2137 1472 2350 1477
rect 2921 1472 2974 1477
rect 593 1467 598 1472
rect 265 1462 310 1467
rect 329 1462 446 1467
rect 521 1462 542 1467
rect 593 1462 622 1467
rect 689 1462 774 1467
rect 841 1462 1006 1467
rect 1177 1462 1486 1467
rect 1569 1462 1718 1467
rect 1737 1462 1846 1467
rect 1945 1462 2062 1467
rect 2089 1462 2158 1467
rect 2361 1462 2614 1467
rect 2713 1462 2742 1467
rect 2913 1462 3230 1467
rect 1025 1457 1158 1462
rect 1737 1457 1742 1462
rect 201 1452 382 1457
rect 433 1452 966 1457
rect 977 1452 1030 1457
rect 1153 1452 1334 1457
rect 1361 1452 1390 1457
rect 1489 1452 1742 1457
rect 1841 1457 1846 1462
rect 2153 1457 2158 1462
rect 2273 1457 2366 1462
rect 1841 1452 1950 1457
rect 1969 1452 2134 1457
rect 2153 1452 2278 1457
rect 2521 1452 2582 1457
rect 2625 1452 2678 1457
rect 2833 1452 2934 1457
rect 2577 1447 2582 1452
rect 73 1442 190 1447
rect 273 1442 358 1447
rect 369 1442 406 1447
rect 417 1442 446 1447
rect 481 1442 582 1447
rect 625 1442 734 1447
rect 849 1442 958 1447
rect 1017 1442 1438 1447
rect 1489 1442 1526 1447
rect 1585 1442 1718 1447
rect 1745 1442 1902 1447
rect 1993 1442 2046 1447
rect 2297 1442 2558 1447
rect 2577 1442 2870 1447
rect 2881 1442 3110 1447
rect 401 1437 406 1442
rect 145 1432 230 1437
rect 401 1432 750 1437
rect 793 1432 846 1437
rect 897 1432 1814 1437
rect 2001 1432 2038 1437
rect 2169 1432 2262 1437
rect 2281 1432 2366 1437
rect 2497 1432 2598 1437
rect 2673 1432 2726 1437
rect 2905 1432 2926 1437
rect 3041 1432 3134 1437
rect 2169 1427 2174 1432
rect 273 1422 302 1427
rect 321 1422 550 1427
rect 561 1422 590 1427
rect 649 1422 678 1427
rect 545 1417 550 1422
rect 65 1412 94 1417
rect 113 1412 166 1417
rect 345 1412 374 1417
rect 385 1412 414 1417
rect 449 1412 534 1417
rect 545 1412 646 1417
rect 65 1397 70 1412
rect 209 1407 326 1412
rect 145 1402 214 1407
rect 321 1402 358 1407
rect 369 1402 374 1412
rect 529 1407 534 1412
rect 673 1407 678 1422
rect 697 1417 702 1427
rect 961 1422 1078 1427
rect 1073 1417 1078 1422
rect 1169 1417 1174 1427
rect 1289 1422 1534 1427
rect 1625 1422 1926 1427
rect 1961 1422 2014 1427
rect 2033 1422 2110 1427
rect 2145 1422 2174 1427
rect 2257 1427 2262 1432
rect 2257 1422 2350 1427
rect 2377 1422 2414 1427
rect 2561 1422 2606 1427
rect 2713 1422 2814 1427
rect 2897 1422 2942 1427
rect 697 1412 710 1417
rect 777 1412 798 1417
rect 905 1412 1054 1417
rect 1073 1412 1174 1417
rect 1249 1412 1278 1417
rect 1297 1412 1654 1417
rect 1865 1412 2310 1417
rect 2337 1412 2374 1417
rect 2625 1412 2734 1417
rect 2753 1412 2886 1417
rect 2953 1412 3110 1417
rect 3257 1412 3358 1417
rect 385 1402 518 1407
rect 529 1402 566 1407
rect 601 1402 630 1407
rect 641 1402 678 1407
rect 705 1407 710 1412
rect 1297 1407 1302 1412
rect 1649 1407 1870 1412
rect 705 1402 774 1407
rect 937 1402 958 1407
rect 1025 1402 1086 1407
rect 1137 1402 1302 1407
rect 1369 1402 1414 1407
rect 1457 1402 1630 1407
rect 1889 1402 1966 1407
rect 1977 1402 2286 1407
rect 2369 1402 2374 1412
rect 2753 1407 2758 1412
rect 2881 1407 2958 1412
rect 2681 1402 2758 1407
rect 1457 1397 1462 1402
rect 2833 1397 2838 1407
rect 3105 1402 3110 1412
rect 3225 1402 3286 1407
rect 65 1392 134 1397
rect 225 1392 310 1397
rect 345 1392 438 1397
rect 449 1392 838 1397
rect 865 1392 1182 1397
rect 1257 1392 1462 1397
rect 1481 1392 1510 1397
rect 1657 1392 1862 1397
rect 1969 1392 2038 1397
rect 2081 1392 2142 1397
rect 2177 1392 2326 1397
rect 2649 1392 2910 1397
rect 3009 1392 3230 1397
rect 129 1387 134 1392
rect 433 1387 438 1392
rect 2345 1387 2438 1392
rect 89 1382 118 1387
rect 129 1382 422 1387
rect 433 1382 470 1387
rect 489 1382 838 1387
rect 937 1382 982 1387
rect 993 1382 1046 1387
rect 1057 1382 1078 1387
rect 1129 1382 1174 1387
rect 1281 1382 1302 1387
rect 1409 1382 1526 1387
rect 1577 1382 1622 1387
rect 1849 1382 2014 1387
rect 2041 1382 2078 1387
rect 2129 1382 2182 1387
rect 2289 1382 2350 1387
rect 2433 1382 2462 1387
rect 2553 1382 2630 1387
rect 2649 1382 2854 1387
rect 417 1377 422 1382
rect 849 1377 942 1382
rect 297 1372 366 1377
rect 417 1372 598 1377
rect 625 1372 774 1377
rect 785 1372 854 1377
rect 961 1372 1046 1377
rect 185 1367 278 1372
rect 769 1367 774 1372
rect 1057 1367 1062 1382
rect 2553 1377 2558 1382
rect 1073 1372 1134 1377
rect 1385 1372 2022 1377
rect 2153 1372 2446 1377
rect 2529 1372 2558 1377
rect 2625 1377 2630 1382
rect 2625 1372 2726 1377
rect 2777 1372 2838 1377
rect 2873 1372 2942 1377
rect 2961 1372 3118 1377
rect 3393 1372 3414 1377
rect 1241 1367 1366 1372
rect 2041 1367 2134 1372
rect 2961 1367 2966 1372
rect 81 1362 150 1367
rect 161 1362 190 1367
rect 273 1362 446 1367
rect 481 1362 534 1367
rect 609 1362 638 1367
rect 673 1362 742 1367
rect 769 1362 950 1367
rect 1009 1362 1062 1367
rect 1081 1362 1102 1367
rect 1113 1362 1246 1367
rect 1361 1362 1486 1367
rect 1505 1362 1662 1367
rect 1769 1362 1798 1367
rect 1873 1362 1974 1367
rect 1993 1362 2046 1367
rect 2129 1362 2614 1367
rect 2865 1362 2966 1367
rect 3113 1367 3118 1372
rect 3113 1362 3142 1367
rect 3289 1362 3398 1367
rect 2609 1357 2742 1362
rect 2865 1357 2870 1362
rect 193 1352 270 1357
rect 289 1352 2246 1357
rect 2257 1352 2286 1357
rect 2393 1352 2590 1357
rect 2737 1352 2870 1357
rect 2953 1352 3062 1357
rect 3097 1352 3262 1357
rect 2241 1347 2246 1352
rect 2281 1347 2398 1352
rect 3409 1347 3414 1372
rect 289 1342 734 1347
rect 849 1342 1286 1347
rect 1313 1342 1366 1347
rect 1385 1342 1574 1347
rect 1585 1342 1646 1347
rect 1665 1342 1702 1347
rect 1745 1342 1854 1347
rect 1881 1342 2174 1347
rect 2241 1342 2262 1347
rect 2417 1342 2534 1347
rect 2697 1342 2718 1347
rect 2889 1342 2942 1347
rect 3001 1342 3174 1347
rect 3393 1342 3414 1347
rect 729 1337 854 1342
rect 2257 1337 2262 1342
rect 161 1332 382 1337
rect 465 1332 510 1337
rect 665 1332 710 1337
rect 873 1332 1118 1337
rect 1225 1332 1694 1337
rect 1721 1332 2070 1337
rect 529 1327 638 1332
rect 2065 1327 2070 1332
rect 2185 1332 2246 1337
rect 2257 1332 2606 1337
rect 3089 1332 3150 1337
rect 3257 1332 3302 1337
rect 2185 1327 2190 1332
rect 81 1322 126 1327
rect 209 1322 238 1327
rect 281 1322 302 1327
rect 385 1322 406 1327
rect 433 1322 534 1327
rect 633 1322 662 1327
rect 673 1322 1678 1327
rect 1761 1322 1838 1327
rect 1889 1322 1998 1327
rect 2065 1322 2190 1327
rect 2329 1322 2438 1327
rect 2553 1322 2614 1327
rect 2729 1322 2774 1327
rect 2849 1322 2918 1327
rect 2929 1322 3038 1327
rect 673 1317 678 1322
rect 1673 1317 1766 1322
rect 361 1312 414 1317
rect 497 1312 550 1317
rect 577 1312 622 1317
rect 657 1312 678 1317
rect 881 1312 982 1317
rect 1009 1312 1270 1317
rect 1281 1312 1406 1317
rect 1425 1312 1446 1317
rect 1489 1312 1654 1317
rect 1785 1312 1862 1317
rect 753 1307 862 1312
rect 1265 1307 1270 1312
rect 1857 1307 1862 1312
rect 1889 1307 1894 1322
rect 3089 1317 3094 1332
rect 3313 1327 3318 1337
rect 3129 1322 3174 1327
rect 3225 1322 3278 1327
rect 3297 1322 3318 1327
rect 3345 1322 3382 1327
rect 1905 1312 2046 1317
rect 2401 1312 2462 1317
rect 2809 1312 2958 1317
rect 3009 1312 3094 1317
rect 3113 1312 3142 1317
rect 3009 1307 3014 1312
rect 121 1302 166 1307
rect 281 1302 310 1307
rect 441 1302 566 1307
rect 609 1302 686 1307
rect 729 1302 758 1307
rect 857 1302 894 1307
rect 913 1302 1254 1307
rect 1265 1302 1550 1307
rect 1673 1302 1814 1307
rect 1857 1302 1926 1307
rect 1953 1302 2086 1307
rect 2161 1302 2302 1307
rect 2417 1302 2470 1307
rect 2625 1302 2750 1307
rect 2769 1302 3014 1307
rect 3041 1302 3174 1307
rect 1569 1297 1678 1302
rect 2161 1297 2166 1302
rect 2625 1297 2630 1302
rect 401 1292 422 1297
rect 465 1292 510 1297
rect 521 1292 678 1297
rect 705 1292 854 1297
rect 993 1292 1046 1297
rect 1121 1292 1166 1297
rect 1193 1292 1326 1297
rect 1385 1292 1574 1297
rect 1793 1292 2022 1297
rect 2073 1292 2166 1297
rect 2353 1292 2462 1297
rect 2601 1292 2630 1297
rect 2745 1297 2750 1302
rect 2745 1292 3142 1297
rect 249 1287 382 1292
rect 225 1282 254 1287
rect 377 1282 590 1287
rect 673 1277 678 1292
rect 873 1287 974 1292
rect 2185 1287 2254 1292
rect 833 1282 878 1287
rect 969 1282 1246 1287
rect 1449 1282 1486 1287
rect 1545 1282 2038 1287
rect 2097 1282 2190 1287
rect 2249 1282 2342 1287
rect 2417 1282 3046 1287
rect 1265 1277 1406 1282
rect 2033 1277 2038 1282
rect 2337 1277 2422 1282
rect 233 1272 630 1277
rect 673 1272 702 1277
rect 809 1272 1110 1277
rect 1121 1272 1270 1277
rect 1401 1272 1430 1277
rect 1489 1272 1526 1277
rect 1569 1272 1670 1277
rect 1681 1272 1750 1277
rect 1849 1272 1878 1277
rect 1889 1272 2022 1277
rect 2033 1272 2238 1277
rect 2609 1272 2806 1277
rect 3065 1272 3094 1277
rect 3225 1272 3334 1277
rect 1105 1267 1110 1272
rect 1489 1267 1494 1272
rect 1681 1267 1686 1272
rect 1745 1267 1854 1272
rect 1873 1267 1878 1272
rect 2017 1267 2022 1272
rect 2801 1267 3070 1272
rect 305 1262 326 1267
rect 361 1262 446 1267
rect 569 1262 678 1267
rect 1001 1262 1078 1267
rect 1105 1262 1494 1267
rect 1505 1262 1686 1267
rect 1873 1262 1942 1267
rect 2017 1262 2230 1267
rect 2305 1262 2542 1267
rect 2561 1262 2782 1267
rect 3113 1262 3206 1267
rect 193 1257 286 1262
rect 673 1257 678 1262
rect 721 1257 886 1262
rect 2537 1257 2542 1262
rect 3113 1257 3118 1262
rect 3201 1257 3310 1262
rect 137 1252 198 1257
rect 281 1252 438 1257
rect 513 1252 542 1257
rect 641 1252 662 1257
rect 673 1252 726 1257
rect 881 1252 1326 1257
rect 1345 1252 1486 1257
rect 1497 1252 1686 1257
rect 1745 1252 1798 1257
rect 1825 1252 2006 1257
rect 2025 1252 2302 1257
rect 2537 1252 2662 1257
rect 2697 1252 2774 1257
rect 2841 1252 2942 1257
rect 2993 1252 3118 1257
rect 3305 1252 3334 1257
rect 561 1247 646 1252
rect 2345 1247 2518 1252
rect 161 1242 326 1247
rect 401 1242 566 1247
rect 665 1242 870 1247
rect 993 1242 1118 1247
rect 1129 1242 1158 1247
rect 1185 1242 1374 1247
rect 1529 1242 1662 1247
rect 1689 1242 2062 1247
rect 1369 1237 1534 1242
rect 1657 1237 1662 1242
rect 2057 1237 2062 1242
rect 2177 1242 2350 1247
rect 2513 1242 2678 1247
rect 2729 1242 2910 1247
rect 3225 1242 3326 1247
rect 2177 1237 2182 1242
rect 2929 1237 3206 1242
rect 217 1232 254 1237
rect 289 1232 310 1237
rect 433 1232 470 1237
rect 529 1232 590 1237
rect 617 1232 750 1237
rect 809 1232 1206 1237
rect 1217 1232 1350 1237
rect 1553 1232 1638 1237
rect 1657 1232 1726 1237
rect 1737 1232 2038 1237
rect 2057 1232 2182 1237
rect 2209 1232 2934 1237
rect 3201 1232 3310 1237
rect 3345 1232 3366 1237
rect 121 1222 230 1227
rect 433 1217 438 1232
rect 1201 1227 1206 1232
rect 449 1222 606 1227
rect 625 1222 670 1227
rect 745 1222 782 1227
rect 793 1222 886 1227
rect 937 1222 1006 1227
rect 1049 1222 1086 1227
rect 1097 1222 1166 1227
rect 1201 1222 1230 1227
rect 1369 1222 1462 1227
rect 1481 1222 1790 1227
rect 1905 1222 1990 1227
rect 2201 1222 2246 1227
rect 2385 1222 2438 1227
rect 2537 1222 2590 1227
rect 2609 1222 2638 1227
rect 2745 1222 2782 1227
rect 2817 1222 2926 1227
rect 2969 1222 3062 1227
rect 3073 1222 3126 1227
rect 3137 1222 3158 1227
rect 3185 1222 3254 1227
rect 3281 1222 3302 1227
rect 3321 1222 3342 1227
rect 1249 1217 1374 1222
rect 1457 1217 1462 1222
rect 2609 1217 2614 1222
rect 73 1207 78 1217
rect 89 1212 150 1217
rect 353 1212 390 1217
rect 433 1212 478 1217
rect 577 1212 710 1217
rect 785 1212 1254 1217
rect 1457 1212 1526 1217
rect 1625 1212 1742 1217
rect 1769 1212 1822 1217
rect 1849 1212 2086 1217
rect 2249 1212 2286 1217
rect 2321 1212 2582 1217
rect 2593 1212 2614 1217
rect 2633 1212 2814 1217
rect 193 1207 262 1212
rect 65 1202 78 1207
rect 137 1202 198 1207
rect 257 1202 286 1207
rect 313 1202 406 1207
rect 65 1197 70 1202
rect 65 1192 94 1197
rect 209 1192 254 1197
rect 297 1192 558 1197
rect 577 1192 582 1212
rect 1521 1207 1630 1212
rect 2105 1207 2230 1212
rect 2833 1207 2918 1212
rect 601 1202 1502 1207
rect 1649 1202 2110 1207
rect 2225 1202 2838 1207
rect 2913 1202 2974 1207
rect 3041 1202 3062 1207
rect 681 1192 758 1197
rect 801 1192 846 1197
rect 881 1192 974 1197
rect 1001 1192 1062 1197
rect 1081 1192 1150 1197
rect 1249 1192 1374 1197
rect 553 1187 558 1192
rect 1145 1187 1254 1192
rect 1369 1187 1374 1192
rect 1505 1192 1638 1197
rect 1825 1192 2270 1197
rect 2393 1192 2750 1197
rect 2785 1192 2830 1197
rect 2881 1192 2902 1197
rect 3081 1192 3126 1197
rect 1505 1187 1510 1192
rect 1633 1187 1638 1192
rect 1737 1187 1830 1192
rect 2265 1187 2398 1192
rect 3153 1187 3158 1222
rect 3201 1212 3230 1217
rect 3201 1207 3206 1212
rect 3201 1202 3278 1207
rect 3297 1197 3302 1222
rect 3361 1217 3366 1232
rect 3337 1212 3366 1217
rect 3369 1202 3398 1207
rect 3233 1192 3366 1197
rect 161 1182 318 1187
rect 329 1182 374 1187
rect 553 1182 1126 1187
rect 1273 1182 1334 1187
rect 1369 1182 1510 1187
rect 1529 1182 1614 1187
rect 1633 1182 1742 1187
rect 1849 1182 1942 1187
rect 1961 1182 2102 1187
rect 2169 1182 2246 1187
rect 2417 1182 2534 1187
rect 2585 1182 3134 1187
rect 3153 1182 3366 1187
rect 1937 1177 1942 1182
rect 49 1172 326 1177
rect 337 1172 366 1177
rect 401 1172 550 1177
rect 561 1172 702 1177
rect 713 1172 766 1177
rect 809 1172 902 1177
rect 1017 1172 1118 1177
rect 1145 1172 1230 1177
rect 1321 1172 1350 1177
rect 1529 1172 1590 1177
rect 1761 1172 1830 1177
rect 1857 1172 1934 1177
rect 1937 1172 2158 1177
rect 2209 1172 2358 1177
rect 2377 1172 2470 1177
rect 2561 1172 2582 1177
rect 2681 1172 2854 1177
rect 2985 1172 3014 1177
rect 49 1157 54 1172
rect 1145 1167 1150 1172
rect 73 1162 126 1167
rect 209 1162 262 1167
rect 337 1162 374 1167
rect 385 1162 1150 1167
rect 1225 1167 1230 1172
rect 1761 1167 1766 1172
rect 1225 1162 1766 1167
rect 1825 1167 1830 1172
rect 1929 1167 1934 1172
rect 3009 1167 3014 1172
rect 3089 1172 3158 1177
rect 3265 1172 3350 1177
rect 3377 1172 3382 1197
rect 3089 1167 3094 1172
rect 3393 1167 3398 1202
rect 1825 1162 1926 1167
rect 1929 1162 2206 1167
rect 2233 1162 2726 1167
rect 2753 1162 2918 1167
rect 3009 1162 3094 1167
rect 3137 1162 3286 1167
rect 3369 1162 3398 1167
rect 209 1157 214 1162
rect 369 1157 374 1162
rect 1921 1157 1926 1162
rect 49 1152 78 1157
rect 145 1152 214 1157
rect 257 1152 350 1157
rect 369 1152 446 1157
rect 513 1152 686 1157
rect 737 1152 990 1157
rect 1097 1152 1334 1157
rect 1777 1152 1910 1157
rect 1921 1152 2174 1157
rect 2185 1152 2358 1157
rect 2513 1152 2590 1157
rect 2633 1152 2798 1157
rect 2809 1152 2958 1157
rect 3113 1152 3254 1157
rect 2377 1147 2494 1152
rect 201 1142 526 1147
rect 617 1142 1326 1147
rect 1521 1142 1550 1147
rect 1769 1142 2382 1147
rect 2489 1142 2790 1147
rect 2801 1142 2894 1147
rect 2905 1142 2942 1147
rect 3033 1142 3214 1147
rect 3337 1142 3358 1147
rect 97 1132 118 1137
rect 209 1132 310 1137
rect 321 1132 350 1137
rect 369 1132 390 1137
rect 433 1132 590 1137
rect 681 1132 750 1137
rect 761 1132 798 1137
rect 897 1132 950 1137
rect 977 1132 1062 1137
rect 1081 1132 1142 1137
rect 1217 1132 1270 1137
rect 1337 1132 1758 1137
rect 1865 1132 2350 1137
rect 2377 1132 2534 1137
rect 2601 1132 2870 1137
rect 2881 1132 2974 1137
rect 3137 1132 3246 1137
rect 113 1127 118 1132
rect 369 1127 374 1132
rect 1753 1127 1870 1132
rect 89 1122 118 1127
rect 249 1122 374 1127
rect 465 1122 582 1127
rect 713 1122 950 1127
rect 1105 1122 1206 1127
rect 1281 1122 1406 1127
rect 1889 1122 2230 1127
rect 2273 1122 2310 1127
rect 2353 1122 2454 1127
rect 2537 1122 2566 1127
rect 2657 1122 2726 1127
rect 2745 1122 2854 1127
rect 3153 1122 3254 1127
rect 601 1117 694 1122
rect 1201 1117 1286 1122
rect 2721 1117 2726 1122
rect 97 1112 126 1117
rect 385 1112 446 1117
rect 577 1112 606 1117
rect 689 1112 1142 1117
rect 1625 1112 1670 1117
rect 1713 1112 1902 1117
rect 2089 1112 2366 1117
rect 2465 1112 2566 1117
rect 2649 1112 2694 1117
rect 2721 1112 2758 1117
rect 2777 1112 3086 1117
rect 3113 1112 3342 1117
rect 2361 1107 2470 1112
rect 2561 1107 2566 1112
rect 2753 1107 2758 1112
rect 353 1102 390 1107
rect 449 1102 566 1107
rect 625 1102 814 1107
rect 857 1102 1118 1107
rect 1217 1102 1246 1107
rect 1449 1102 1606 1107
rect 2001 1102 2070 1107
rect 2097 1102 2342 1107
rect 2561 1102 2614 1107
rect 2681 1102 2726 1107
rect 2753 1102 2782 1107
rect 2801 1102 2894 1107
rect 3017 1102 3086 1107
rect 3145 1102 3190 1107
rect 1449 1097 1454 1102
rect 1601 1097 1846 1102
rect 2337 1097 2342 1102
rect 2609 1097 2614 1102
rect 401 1092 422 1097
rect 433 1092 486 1097
rect 513 1092 886 1097
rect 921 1092 1030 1097
rect 1041 1092 1102 1097
rect 1289 1092 1406 1097
rect 1425 1092 1454 1097
rect 1841 1092 2038 1097
rect 2057 1092 2102 1097
rect 2121 1092 2254 1097
rect 2337 1092 2438 1097
rect 2457 1092 2590 1097
rect 2609 1092 2822 1097
rect 2841 1092 2918 1097
rect 3113 1092 3222 1097
rect 1025 1087 1030 1092
rect 1289 1087 1294 1092
rect 209 1082 278 1087
rect 393 1082 454 1087
rect 465 1082 606 1087
rect 665 1082 726 1087
rect 777 1082 894 1087
rect 937 1082 1014 1087
rect 1025 1082 1134 1087
rect 1193 1082 1294 1087
rect 1401 1087 1406 1092
rect 1473 1087 1582 1092
rect 2033 1087 2038 1092
rect 2433 1087 2438 1092
rect 1401 1082 1478 1087
rect 1577 1082 1830 1087
rect 2033 1082 2326 1087
rect 2433 1082 2662 1087
rect 2673 1082 2750 1087
rect 2777 1082 2822 1087
rect 2929 1082 3014 1087
rect 3129 1082 3182 1087
rect 209 1077 214 1082
rect 137 1072 214 1077
rect 273 1077 278 1082
rect 465 1077 470 1082
rect 1825 1077 2014 1082
rect 2817 1077 2934 1082
rect 273 1072 470 1077
rect 481 1072 782 1077
rect 801 1072 1814 1077
rect 2009 1072 2086 1077
rect 2097 1072 2158 1077
rect 2193 1072 2222 1077
rect 2281 1072 2526 1077
rect 2545 1072 2798 1077
rect 3129 1072 3206 1077
rect 2097 1067 2102 1072
rect 2545 1067 2550 1072
rect 353 1062 518 1067
rect 537 1062 742 1067
rect 753 1062 846 1067
rect 881 1062 910 1067
rect 945 1062 966 1067
rect 1025 1062 1046 1067
rect 1113 1062 1142 1067
rect 1185 1062 1230 1067
rect 1537 1062 1606 1067
rect 1681 1062 2102 1067
rect 2329 1062 2550 1067
rect 2601 1062 2630 1067
rect 2673 1062 2758 1067
rect 2817 1062 2910 1067
rect 753 1057 758 1062
rect 1249 1057 1358 1062
rect 1393 1057 1470 1062
rect 1681 1057 1686 1062
rect 2121 1057 2310 1062
rect 2817 1057 2822 1062
rect 225 1052 262 1057
rect 465 1052 654 1057
rect 689 1052 758 1057
rect 801 1052 878 1057
rect 913 1052 1054 1057
rect 1129 1052 1254 1057
rect 1353 1052 1398 1057
rect 1465 1052 1526 1057
rect 1585 1052 1686 1057
rect 1769 1052 2126 1057
rect 2305 1052 2822 1057
rect 2905 1057 2910 1062
rect 2905 1052 2934 1057
rect 2969 1052 3094 1057
rect 3169 1052 3270 1057
rect 289 1047 358 1052
rect 1521 1047 1590 1052
rect 2969 1047 2974 1052
rect 265 1042 294 1047
rect 353 1042 1342 1047
rect 1409 1042 1454 1047
rect 1609 1042 2894 1047
rect 2945 1042 2974 1047
rect 289 1032 342 1037
rect 457 1032 598 1037
rect 697 1032 734 1037
rect 745 1032 926 1037
rect 969 1032 2214 1037
rect 2225 1032 2390 1037
rect 2465 1032 2702 1037
rect 2761 1032 2798 1037
rect 2945 1032 3070 1037
rect 289 1017 294 1032
rect 2225 1027 2230 1032
rect 3089 1027 3094 1052
rect 3105 1042 3222 1047
rect 3177 1032 3302 1037
rect 3177 1027 3182 1032
rect 305 1022 534 1027
rect 577 1022 646 1027
rect 705 1022 894 1027
rect 945 1022 1022 1027
rect 1049 1022 1070 1027
rect 1097 1022 1222 1027
rect 1233 1022 1278 1027
rect 1297 1022 1510 1027
rect 1577 1022 1822 1027
rect 1905 1022 1934 1027
rect 2001 1022 2230 1027
rect 2265 1022 2294 1027
rect 2521 1022 2814 1027
rect 2841 1022 2958 1027
rect 3089 1022 3182 1027
rect 945 1017 950 1022
rect 177 1012 214 1017
rect 289 1012 358 1017
rect 417 1012 950 1017
rect 993 1017 998 1022
rect 1297 1017 1302 1022
rect 1817 1017 1910 1022
rect 2289 1017 2454 1022
rect 2521 1017 2526 1022
rect 993 1012 1302 1017
rect 1409 1012 1486 1017
rect 1553 1012 1798 1017
rect 1945 1012 2062 1017
rect 2073 1012 2238 1017
rect 2449 1012 2526 1017
rect 2593 1012 2686 1017
rect 2873 1012 2966 1017
rect 2993 1012 3054 1017
rect 113 1002 222 1007
rect 281 1002 326 1007
rect 353 997 358 1012
rect 1329 1007 1414 1012
rect 425 1002 486 1007
rect 521 1002 694 1007
rect 737 1002 854 1007
rect 905 1002 1334 1007
rect 1433 1002 1870 1007
rect 1905 1002 2166 1007
rect 2249 1002 2414 1007
rect 2545 1002 2614 1007
rect 2825 1002 3006 1007
rect 3153 1002 3230 1007
rect 193 992 334 997
rect 353 992 390 997
rect 569 992 646 997
rect 737 987 742 1002
rect 2161 997 2254 1002
rect 3393 997 3398 1017
rect 777 992 950 997
rect 1017 992 1054 997
rect 1065 992 1342 997
rect 1361 992 1398 997
rect 1545 992 1646 997
rect 1793 992 1966 997
rect 2001 992 2070 997
rect 2105 992 2142 997
rect 2393 992 3022 997
rect 3049 992 3118 997
rect 3297 992 3398 997
rect 1361 987 1366 992
rect 1417 987 1526 992
rect 1665 987 1758 992
rect 3049 987 3054 992
rect 289 982 318 987
rect 313 977 318 982
rect 401 982 590 987
rect 697 982 742 987
rect 969 982 1014 987
rect 1057 982 1126 987
rect 1297 982 1366 987
rect 1377 982 1422 987
rect 1521 982 1670 987
rect 1753 982 1782 987
rect 1793 982 2246 987
rect 2257 982 2326 987
rect 2577 982 2630 987
rect 2729 982 2782 987
rect 2809 982 2838 987
rect 3033 982 3054 987
rect 3113 987 3118 992
rect 3113 982 3142 987
rect 3337 982 3366 987
rect 401 977 406 982
rect 761 977 950 982
rect 1145 977 1262 982
rect 2241 977 2246 982
rect 2345 977 2558 982
rect 2833 977 2950 982
rect 3033 977 3038 982
rect 313 972 406 977
rect 537 972 766 977
rect 945 972 1150 977
rect 1257 972 1502 977
rect 1521 972 1606 977
rect 1625 972 1750 977
rect 1833 972 2182 977
rect 2241 972 2350 977
rect 2553 972 2678 977
rect 2945 972 3038 977
rect 3065 972 3206 977
rect 569 962 598 967
rect 609 962 1134 967
rect 1185 962 1614 967
rect 1665 962 1822 967
rect 1833 962 1862 967
rect 1985 962 2030 967
rect 2057 962 2102 967
rect 2113 962 2174 967
rect 2329 962 2462 967
rect 2481 962 2518 967
rect 2537 962 2606 967
rect 2641 962 2710 967
rect 2745 962 2790 967
rect 2841 962 2926 967
rect 2193 957 2310 962
rect 2841 957 2846 962
rect 161 952 342 957
rect 377 952 526 957
rect 545 952 670 957
rect 697 952 718 957
rect 801 952 1094 957
rect 1249 952 1494 957
rect 1529 952 2198 957
rect 2305 952 2710 957
rect 2793 952 2846 957
rect 2921 957 2926 962
rect 3153 957 3230 962
rect 2921 952 2950 957
rect 3097 952 3158 957
rect 3225 952 3254 957
rect 1089 947 1254 952
rect 2705 947 2798 952
rect 97 942 134 947
rect 465 942 838 947
rect 833 937 838 942
rect 905 942 1070 947
rect 1345 942 1582 947
rect 1625 942 1686 947
rect 1697 942 2206 947
rect 2217 942 2422 947
rect 2465 942 2542 947
rect 2569 942 2662 947
rect 2833 942 2982 947
rect 3169 942 3198 947
rect 3329 942 3358 947
rect 905 937 910 942
rect 233 932 430 937
rect 497 932 622 937
rect 657 932 702 937
rect 785 932 814 937
rect 833 932 910 937
rect 945 932 982 937
rect 1097 932 1118 937
rect 1233 932 1302 937
rect 1545 932 1670 937
rect 697 927 790 932
rect 1377 927 1526 932
rect 1697 927 1702 942
rect 1737 932 1894 937
rect 1929 932 2510 937
rect 2529 932 2582 937
rect 2721 932 2750 937
rect 2801 932 2934 937
rect 3049 932 3198 937
rect 3233 932 3310 937
rect 3233 927 3238 932
rect 185 922 222 927
rect 249 922 294 927
rect 337 922 398 927
rect 457 922 534 927
rect 1129 922 1382 927
rect 1521 922 1702 927
rect 1825 922 1926 927
rect 2081 922 2150 927
rect 2185 922 2630 927
rect 2777 922 2886 927
rect 2897 922 3038 927
rect 3209 922 3238 927
rect 3305 927 3310 932
rect 3305 922 3374 927
rect 257 912 278 917
rect 105 902 238 907
rect 193 892 262 897
rect 273 887 278 912
rect 233 882 278 887
rect 289 887 294 922
rect 553 917 678 922
rect 1041 917 1134 922
rect 1945 917 2062 922
rect 2649 917 2758 922
rect 2897 917 2902 922
rect 3033 917 3214 922
rect 433 912 558 917
rect 673 912 702 917
rect 721 912 846 917
rect 977 912 1022 917
rect 1041 907 1046 917
rect 1177 912 1246 917
rect 1393 912 1950 917
rect 2057 912 2654 917
rect 2753 912 2902 917
rect 3249 912 3294 917
rect 425 902 574 907
rect 585 902 1046 907
rect 1057 902 1110 907
rect 1129 902 1214 907
rect 1233 902 1366 907
rect 1377 902 1526 907
rect 1545 902 1574 907
rect 1633 902 1710 907
rect 1793 902 1822 907
rect 1937 902 2078 907
rect 2129 902 2158 907
rect 2217 902 2438 907
rect 2521 902 2582 907
rect 2633 902 2710 907
rect 2737 902 2774 907
rect 2849 902 2886 907
rect 2921 902 3062 907
rect 3105 902 3190 907
rect 3209 902 3358 907
rect 2921 897 2926 902
rect 377 892 430 897
rect 441 892 534 897
rect 593 892 878 897
rect 977 892 1006 897
rect 1017 892 1142 897
rect 1193 892 1430 897
rect 1609 892 2390 897
rect 2409 892 2662 897
rect 2769 892 2862 897
rect 2889 892 2926 897
rect 3057 897 3062 902
rect 3057 892 3086 897
rect 3217 892 3262 897
rect 1449 887 1590 892
rect 289 882 422 887
rect 577 882 1254 887
rect 1297 882 1454 887
rect 1585 882 3206 887
rect 441 877 510 882
rect 177 872 270 877
rect 313 872 446 877
rect 505 872 1750 877
rect 1969 872 2190 877
rect 2281 872 2534 877
rect 2577 872 2886 877
rect 3041 872 3238 877
rect 1745 867 1974 872
rect 2185 867 2286 872
rect 2529 867 2534 872
rect 257 862 334 867
rect 441 862 494 867
rect 569 862 630 867
rect 673 862 886 867
rect 961 862 1014 867
rect 1065 862 1086 867
rect 1129 862 1222 867
rect 1241 862 1278 867
rect 1337 862 1374 867
rect 1409 862 1726 867
rect 1993 862 2166 867
rect 2305 862 2398 867
rect 2409 862 2510 867
rect 2529 862 2622 867
rect 2825 862 3174 867
rect 3249 862 3406 867
rect 673 857 678 862
rect 3169 857 3254 862
rect 161 852 238 857
rect 257 852 286 857
rect 609 852 678 857
rect 689 852 1406 857
rect 1497 852 1774 857
rect 1873 852 1990 857
rect 2041 852 2070 857
rect 2081 852 2110 857
rect 2145 852 2422 857
rect 2433 852 2494 857
rect 2585 852 2654 857
rect 2809 852 2934 857
rect 3049 852 3150 857
rect 161 847 166 852
rect 129 842 166 847
rect 233 847 238 852
rect 233 842 286 847
rect 305 842 398 847
rect 497 842 702 847
rect 713 842 894 847
rect 929 842 1022 847
rect 1057 842 1198 847
rect 1273 842 1582 847
rect 1817 842 2230 847
rect 2321 842 2342 847
rect 2353 842 2550 847
rect 2641 842 3182 847
rect 1057 837 1062 842
rect 1601 837 1782 842
rect 177 832 334 837
rect 361 832 630 837
rect 681 832 726 837
rect 737 832 806 837
rect 833 832 1062 837
rect 1073 832 1142 837
rect 1249 832 1286 837
rect 1321 832 1390 837
rect 1505 832 1606 837
rect 1777 832 1806 837
rect 833 827 838 832
rect 1385 827 1510 832
rect 1801 827 1806 832
rect 1937 832 2310 837
rect 2441 832 2686 837
rect 1937 827 1942 832
rect 2681 827 2686 832
rect 2785 832 2878 837
rect 2961 832 3022 837
rect 3041 832 3102 837
rect 3113 832 3222 837
rect 2785 827 2790 832
rect 193 822 214 827
rect 401 822 462 827
rect 521 822 838 827
rect 857 822 966 827
rect 1057 822 1366 827
rect 1529 822 1742 827
rect 1801 822 1942 827
rect 1961 822 2046 827
rect 2097 822 2150 827
rect 2281 822 2326 827
rect 2361 822 2470 827
rect 2553 822 2614 827
rect 2681 822 2790 827
rect 2849 822 2958 827
rect 2169 817 2262 822
rect 2849 817 2854 822
rect 265 812 310 817
rect 441 812 518 817
rect 553 812 598 817
rect 721 812 782 817
rect 817 812 1302 817
rect 1385 812 1542 817
rect 1553 812 1646 817
rect 2009 812 2054 817
rect 2137 812 2174 817
rect 2257 812 2542 817
rect 2809 812 2854 817
rect 817 807 822 812
rect 1297 807 1302 812
rect 1537 807 1542 812
rect 2049 807 2142 812
rect 2537 807 2662 812
rect 209 802 246 807
rect 281 802 326 807
rect 577 802 822 807
rect 841 802 1286 807
rect 1297 802 1430 807
rect 1537 802 1654 807
rect 1793 802 2030 807
rect 2161 802 2518 807
rect 2657 802 2726 807
rect 2737 802 2774 807
rect 2889 802 2950 807
rect 3009 802 3014 827
rect 3105 822 3134 827
rect 3313 822 3366 827
rect 3313 817 3318 822
rect 3025 812 3070 817
rect 401 797 558 802
rect 2737 797 2742 802
rect 3025 797 3030 812
rect 3153 807 3158 817
rect 3249 812 3318 817
rect 3145 802 3158 807
rect 3281 802 3398 807
rect 185 792 238 797
rect 265 792 406 797
rect 553 792 862 797
rect 897 792 1022 797
rect 1129 792 1326 797
rect 1441 792 1526 797
rect 1537 792 1606 797
rect 2041 792 2070 797
rect 2137 792 2222 797
rect 2321 792 2366 797
rect 2537 792 2742 797
rect 2977 792 3006 797
rect 3017 792 3030 797
rect 3049 792 3110 797
rect 3129 792 3174 797
rect 3289 792 3342 797
rect 1321 787 1446 792
rect 2385 787 2518 792
rect 105 782 182 787
rect 193 782 238 787
rect 297 782 358 787
rect 433 782 726 787
rect 825 782 950 787
rect 985 782 1054 787
rect 1065 782 1118 787
rect 1249 782 1302 787
rect 1465 782 1686 787
rect 1721 782 1822 787
rect 1929 782 2278 787
rect 2289 782 2390 787
rect 2513 782 2670 787
rect 2761 782 2854 787
rect 3017 782 3022 792
rect 3049 782 3198 787
rect 3321 782 3366 787
rect 2761 777 2766 782
rect 129 772 254 777
rect 297 772 334 777
rect 409 772 438 777
rect 497 772 582 777
rect 633 772 1006 777
rect 1137 772 1438 777
rect 1465 772 1494 777
rect 1521 772 1710 777
rect 1721 772 1790 777
rect 1801 772 1822 777
rect 1993 772 2230 777
rect 2241 772 2294 777
rect 2329 772 2414 777
rect 2433 772 2766 777
rect 2849 777 2854 782
rect 2849 772 3030 777
rect 2289 767 2294 772
rect 73 762 1342 767
rect 1481 762 2262 767
rect 2289 762 2622 767
rect 2777 762 2838 767
rect 3025 762 3046 767
rect 3113 762 3214 767
rect 3265 762 3318 767
rect 2617 757 2782 762
rect 3113 757 3118 762
rect 97 752 134 757
rect 177 752 622 757
rect 753 752 998 757
rect 1153 752 1222 757
rect 1313 752 1582 757
rect 1681 752 1766 757
rect 1977 752 2166 757
rect 2209 752 2358 757
rect 2369 752 2438 757
rect 2553 752 2582 757
rect 2929 752 2982 757
rect 3009 752 3078 757
rect 3089 752 3118 757
rect 3209 757 3214 762
rect 3209 752 3302 757
rect 641 747 734 752
rect 1017 747 1134 752
rect 1577 747 1670 752
rect 2465 747 2558 752
rect 113 742 190 747
rect 217 742 502 747
rect 609 742 646 747
rect 729 742 774 747
rect 833 742 1022 747
rect 1129 742 1558 747
rect 1665 742 1726 747
rect 1849 742 2470 747
rect 2649 742 2782 747
rect 2841 742 2966 747
rect 65 722 102 727
rect 113 722 118 742
rect 3009 737 3014 752
rect 3081 742 3110 747
rect 177 732 318 737
rect 505 732 678 737
rect 729 732 1302 737
rect 1489 732 1702 737
rect 1761 732 2326 737
rect 2369 732 2398 737
rect 2481 732 3014 737
rect 3105 737 3110 742
rect 3169 742 3198 747
rect 3169 737 3174 742
rect 3105 732 3174 737
rect 337 727 462 732
rect 1297 727 1302 732
rect 1361 727 1470 732
rect 2481 727 2486 732
rect 145 722 342 727
rect 457 722 1278 727
rect 1297 722 1366 727
rect 1465 722 1518 727
rect 1569 722 2486 727
rect 2865 722 3006 727
rect 3265 722 3310 727
rect 2489 717 2870 722
rect 161 712 198 717
rect 321 712 382 717
rect 321 707 326 712
rect 401 707 406 717
rect 417 712 446 717
rect 561 712 1222 717
rect 1377 712 1814 717
rect 441 707 566 712
rect 1809 707 1814 712
rect 1913 712 2494 717
rect 2889 712 2950 717
rect 1913 707 1918 712
rect 65 702 214 707
rect 281 702 326 707
rect 377 702 406 707
rect 585 702 614 707
rect 705 702 734 707
rect 761 702 798 707
rect 857 702 902 707
rect 969 702 990 707
rect 1017 702 1534 707
rect 1617 702 1790 707
rect 1809 702 1918 707
rect 1953 702 2102 707
rect 2121 702 2182 707
rect 2257 702 2518 707
rect 2561 702 2830 707
rect 3153 702 3302 707
rect 609 697 710 702
rect 2513 697 2518 702
rect 89 692 182 697
rect 217 692 246 697
rect 297 692 326 697
rect 321 687 326 692
rect 409 692 518 697
rect 945 692 1102 697
rect 1129 692 1270 697
rect 1409 692 1438 697
rect 1545 692 1574 697
rect 1649 692 1750 697
rect 1937 692 2246 697
rect 2513 692 2534 697
rect 2793 692 2862 697
rect 409 687 414 692
rect 1289 687 1382 692
rect 1433 687 1550 692
rect 2329 687 2454 692
rect 2857 687 2862 692
rect 2961 692 3102 697
rect 2961 687 2966 692
rect 137 682 166 687
rect 161 677 166 682
rect 233 682 262 687
rect 321 682 414 687
rect 537 682 734 687
rect 801 682 846 687
rect 977 682 1294 687
rect 1377 682 1406 687
rect 1569 682 2158 687
rect 2305 682 2334 687
rect 2449 682 2838 687
rect 2857 682 2966 687
rect 233 677 238 682
rect 537 677 542 682
rect 161 672 238 677
rect 433 672 542 677
rect 729 677 734 682
rect 1569 677 1574 682
rect 729 672 758 677
rect 897 672 958 677
rect 1001 672 1574 677
rect 1585 672 1670 677
rect 1705 672 1766 677
rect 2225 672 2438 677
rect 2529 672 2558 677
rect 1785 667 2190 672
rect 2433 667 2534 672
rect 489 662 1254 667
rect 1345 662 1374 667
rect 1553 662 1790 667
rect 2185 662 2414 667
rect 2657 662 2734 667
rect 1249 657 1350 662
rect 2657 657 2662 662
rect 129 652 262 657
rect 305 652 366 657
rect 385 652 478 657
rect 649 652 670 657
rect 881 652 1118 657
rect 1169 652 1230 657
rect 1481 652 1542 657
rect 1561 652 1646 657
rect 1665 652 1814 657
rect 1841 652 2174 657
rect 2297 652 2502 657
rect 2521 652 2614 657
rect 2633 652 2662 657
rect 2729 657 2734 662
rect 2729 652 2910 657
rect 2929 652 3046 657
rect 449 647 454 652
rect 497 647 630 652
rect 689 647 758 652
rect 1665 647 1670 652
rect 2521 647 2526 652
rect 137 642 222 647
rect 401 642 422 647
rect 449 642 502 647
rect 625 642 694 647
rect 753 642 822 647
rect 929 642 1326 647
rect 1361 642 1670 647
rect 1721 642 1822 647
rect 1833 642 2062 647
rect 2129 642 2326 647
rect 2393 642 2526 647
rect 2609 647 2614 652
rect 2929 647 2934 652
rect 2609 642 2814 647
rect 2905 642 2934 647
rect 3041 647 3046 652
rect 3041 642 3190 647
rect 113 632 310 637
rect 345 632 574 637
rect 617 632 742 637
rect 833 632 1958 637
rect 2009 632 2590 637
rect 2681 632 3030 637
rect 737 627 838 632
rect 2585 627 2686 632
rect 3073 627 3174 632
rect 153 622 462 627
rect 561 622 718 627
rect 873 622 1038 627
rect 1089 622 1150 627
rect 1265 622 1358 627
rect 1497 622 1614 627
rect 1649 622 1718 627
rect 1793 622 1878 627
rect 1929 622 2046 627
rect 2089 622 2206 627
rect 2353 622 2494 627
rect 2841 622 2958 627
rect 3049 622 3078 627
rect 3169 622 3198 627
rect 3233 622 3342 627
rect 1145 617 1270 622
rect 1353 617 1502 622
rect 2225 617 2334 622
rect 3049 617 3054 622
rect 185 612 230 617
rect 369 612 486 617
rect 617 612 678 617
rect 777 612 958 617
rect 1065 612 1126 617
rect 1289 612 1334 617
rect 1521 612 2230 617
rect 2329 612 3054 617
rect 3193 617 3198 622
rect 3193 612 3358 617
rect 369 607 374 612
rect 1521 607 1526 612
rect 209 602 278 607
rect 305 602 374 607
rect 433 602 454 607
rect 497 602 550 607
rect 761 602 854 607
rect 961 602 1046 607
rect 1185 602 1230 607
rect 1345 602 1526 607
rect 1545 602 1774 607
rect 1785 602 1870 607
rect 1921 602 2470 607
rect 2513 602 2638 607
rect 2785 602 2894 607
rect 2969 602 3182 607
rect 305 597 310 602
rect 545 597 550 602
rect 2657 597 2766 602
rect 225 592 310 597
rect 345 592 534 597
rect 545 592 790 597
rect 809 592 1406 597
rect 1505 592 1998 597
rect 2017 592 2238 597
rect 2257 592 2662 597
rect 2761 592 3158 597
rect 785 587 790 592
rect 1401 587 1510 592
rect 417 582 446 587
rect 537 582 566 587
rect 785 582 878 587
rect 985 582 1102 587
rect 1225 582 1382 587
rect 1529 582 2310 587
rect 2369 582 2422 587
rect 2441 582 2958 587
rect 441 577 542 582
rect 2369 577 2374 582
rect 273 572 390 577
rect 385 567 390 572
rect 585 572 702 577
rect 721 572 846 577
rect 993 572 1046 577
rect 1177 572 1518 577
rect 1609 572 2030 577
rect 2297 572 2374 577
rect 2393 572 2558 577
rect 2673 572 2878 577
rect 2953 572 3198 577
rect 3313 572 3358 577
rect 585 567 590 572
rect 313 562 366 567
rect 385 562 590 567
rect 697 567 702 572
rect 1065 567 1158 572
rect 1513 567 1614 572
rect 2049 567 2278 572
rect 697 562 1070 567
rect 1153 562 1366 567
rect 1633 562 1958 567
rect 2009 562 2054 567
rect 2273 562 2654 567
rect 2721 562 2982 567
rect 3153 557 3238 562
rect 161 552 310 557
rect 585 552 1454 557
rect 1473 552 1614 557
rect 1681 552 2750 557
rect 3129 552 3158 557
rect 3233 552 3310 557
rect 1473 547 1478 552
rect 129 542 214 547
rect 297 542 414 547
rect 625 542 686 547
rect 753 542 1254 547
rect 1329 542 1478 547
rect 1609 547 1614 552
rect 1609 542 1998 547
rect 2161 542 2230 547
rect 2281 542 2310 547
rect 2353 542 2510 547
rect 2521 542 2630 547
rect 2833 542 2990 547
rect 3065 542 3094 547
rect 3153 542 3222 547
rect 1249 537 1254 542
rect 2017 537 2142 542
rect 489 532 718 537
rect 785 532 830 537
rect 841 532 1022 537
rect 1113 532 1238 537
rect 1249 532 1598 537
rect 1697 532 2022 537
rect 2137 532 2518 537
rect 3001 532 3062 537
rect 785 527 790 532
rect 1017 527 1118 532
rect 1233 527 1238 532
rect 313 522 374 527
rect 593 522 654 527
rect 737 522 790 527
rect 809 522 854 527
rect 929 522 998 527
rect 1137 522 1206 527
rect 1233 522 1302 527
rect 1313 522 1342 527
rect 1433 522 1478 527
rect 1529 522 1830 527
rect 1841 522 1918 527
rect 1929 522 2334 527
rect 2449 522 2630 527
rect 3217 522 3294 527
rect 73 512 126 517
rect 145 512 214 517
rect 305 512 326 517
rect 825 512 894 517
rect 961 512 966 522
rect 1337 517 1438 522
rect 977 512 1062 517
rect 1113 512 1246 517
rect 1569 512 1790 517
rect 513 507 646 512
rect 1569 507 1574 512
rect 265 502 518 507
rect 641 502 670 507
rect 705 502 1006 507
rect 1017 502 1166 507
rect 1265 502 1406 507
rect 1265 497 1270 502
rect 105 492 134 497
rect 129 487 134 492
rect 273 492 342 497
rect 529 492 814 497
rect 937 492 1270 497
rect 1401 497 1406 502
rect 1457 502 1574 507
rect 1825 507 1830 522
rect 2449 517 2454 522
rect 1849 512 2046 517
rect 2097 512 2454 517
rect 2545 512 2646 517
rect 2665 512 2758 517
rect 2777 512 2910 517
rect 2929 512 2974 517
rect 3081 512 3198 517
rect 2777 507 2782 512
rect 1825 502 1870 507
rect 1897 502 2398 507
rect 2745 502 2782 507
rect 2905 507 2910 512
rect 3081 507 3086 512
rect 2905 502 3086 507
rect 3193 507 3198 512
rect 3193 502 3262 507
rect 3289 502 3326 507
rect 1457 497 1462 502
rect 1657 497 1806 502
rect 1401 492 1462 497
rect 1593 492 1662 497
rect 1801 492 2102 497
rect 2145 492 2174 497
rect 2225 492 2486 497
rect 2537 492 2870 497
rect 3201 492 3382 497
rect 273 487 278 492
rect 2889 487 3118 492
rect 129 482 278 487
rect 561 482 646 487
rect 753 482 1174 487
rect 1281 482 1390 487
rect 1473 482 1582 487
rect 1673 482 2030 487
rect 2161 482 2422 487
rect 2441 482 2566 487
rect 2769 482 2894 487
rect 3113 482 3190 487
rect 1169 477 1286 482
rect 1385 477 1478 482
rect 2081 477 2166 482
rect 2417 477 2422 482
rect 3185 477 3190 482
rect 3329 482 3390 487
rect 3329 477 3334 482
rect 897 472 990 477
rect 1121 472 1150 477
rect 1641 472 1966 477
rect 2017 472 2086 477
rect 2281 472 2342 477
rect 2417 472 2798 477
rect 1009 467 1126 472
rect 2017 467 2022 472
rect 2793 467 2798 472
rect 2897 472 3102 477
rect 3185 472 3334 477
rect 3353 472 3374 477
rect 2897 467 2902 472
rect 377 462 1014 467
rect 1169 462 1614 467
rect 1633 462 2022 467
rect 2033 462 2270 467
rect 2353 462 2774 467
rect 2793 462 2902 467
rect 2993 462 3022 467
rect 1169 457 1174 462
rect 833 452 1174 457
rect 1609 457 1614 462
rect 2265 457 2358 462
rect 1609 452 1726 457
rect 1817 452 2094 457
rect 2473 452 2726 457
rect 697 442 774 447
rect 833 437 838 452
rect 1481 447 1590 452
rect 1721 447 1822 452
rect 2769 447 2774 462
rect 2993 457 2998 462
rect 2921 452 2998 457
rect 3137 452 3230 457
rect 2921 447 2926 452
rect 857 442 1006 447
rect 1041 442 1110 447
rect 1185 442 1486 447
rect 1585 442 1702 447
rect 1841 442 2270 447
rect 2369 442 2750 447
rect 2769 442 2926 447
rect 3105 442 3198 447
rect 1105 437 1190 442
rect 2369 437 2374 442
rect 193 432 238 437
rect 377 432 406 437
rect 537 432 678 437
rect 705 432 838 437
rect 849 432 878 437
rect 945 432 982 437
rect 993 432 1086 437
rect 1337 432 1366 437
rect 1497 432 1526 437
rect 1577 432 2110 437
rect 2201 432 2374 437
rect 2409 432 2534 437
rect 2625 432 2702 437
rect 2945 432 3006 437
rect 3017 432 3062 437
rect 3097 432 3214 437
rect 537 427 542 432
rect 89 422 262 427
rect 513 422 542 427
rect 673 427 678 432
rect 1361 427 1502 432
rect 3057 427 3062 432
rect 673 422 790 427
rect 889 422 1334 427
rect 1593 422 1710 427
rect 1737 422 1766 427
rect 1897 422 1926 427
rect 2041 422 2134 427
rect 2233 422 2262 427
rect 2473 422 2526 427
rect 2953 422 3046 427
rect 3057 422 3126 427
rect 3177 422 3230 427
rect 1761 417 1902 422
rect 2257 417 2478 422
rect 97 412 166 417
rect 369 412 446 417
rect 481 412 550 417
rect 857 412 878 417
rect 1353 412 1574 417
rect 2497 412 2566 417
rect 2905 412 3070 417
rect 569 407 750 412
rect 1009 407 1358 412
rect 1569 407 1574 412
rect 1993 407 2102 412
rect 329 402 574 407
rect 745 402 1014 407
rect 1569 402 1998 407
rect 2097 402 2374 407
rect 2585 402 2774 407
rect 3145 402 3214 407
rect 1377 397 1550 402
rect 2465 397 2590 402
rect 2769 397 2774 402
rect 3025 397 3102 402
rect 201 392 262 397
rect 305 392 454 397
rect 537 392 598 397
rect 625 392 734 397
rect 841 392 894 397
rect 1025 392 1382 397
rect 1545 392 1582 397
rect 2009 392 2086 397
rect 2177 392 2206 397
rect 2345 392 2470 397
rect 2769 392 3030 397
rect 3097 392 3254 397
rect 449 387 542 392
rect 913 387 1006 392
rect 2081 387 2182 392
rect 3249 387 3254 392
rect 361 382 430 387
rect 561 382 918 387
rect 1001 382 1046 387
rect 1065 382 1766 387
rect 1841 382 1974 387
rect 1985 382 2062 387
rect 2481 382 2574 387
rect 2609 382 2758 387
rect 2833 382 2862 387
rect 3041 382 3086 387
rect 3113 382 3142 387
rect 1041 377 1046 382
rect 2753 377 2838 382
rect 3137 377 3142 382
rect 3209 382 3238 387
rect 3249 382 3318 387
rect 3209 377 3214 382
rect 433 372 1022 377
rect 1041 372 1086 377
rect 1121 372 1254 377
rect 1305 372 1526 377
rect 1913 372 2118 377
rect 2129 372 2238 377
rect 2273 372 2334 377
rect 3137 372 3214 377
rect 1521 367 1894 372
rect 2273 367 2278 372
rect 2601 367 2694 372
rect 153 362 350 367
rect 425 362 702 367
rect 849 362 1142 367
rect 1233 362 1502 367
rect 1889 362 2142 367
rect 2177 362 2278 367
rect 2297 362 2430 367
rect 2577 362 2606 367
rect 2689 362 2814 367
rect 2881 362 2950 367
rect 721 357 830 362
rect 1137 357 1222 362
rect 2881 357 2886 362
rect 209 352 286 357
rect 353 352 534 357
rect 625 352 726 357
rect 825 352 982 357
rect 1065 352 1118 357
rect 1217 352 1510 357
rect 1521 352 1574 357
rect 1657 352 2678 357
rect 2769 352 2886 357
rect 2945 357 2950 362
rect 2945 352 2974 357
rect 3041 352 3406 357
rect 2673 347 2774 352
rect 121 342 1062 347
rect 1129 342 1478 347
rect 1817 342 1934 347
rect 2009 342 2078 347
rect 2185 342 2294 347
rect 2385 342 2462 347
rect 2553 342 2654 347
rect 2793 342 2894 347
rect 3337 342 3382 347
rect 1057 337 1134 342
rect 1601 337 1694 342
rect 1729 337 1798 342
rect 193 332 222 337
rect 361 332 526 337
rect 633 332 1038 337
rect 1177 332 1342 337
rect 1577 332 1606 337
rect 1689 332 1734 337
rect 1793 332 3118 337
rect 3129 332 3174 337
rect 3193 332 3318 337
rect 217 327 366 332
rect 1361 327 1558 332
rect 3193 327 3198 332
rect 129 322 198 327
rect 385 322 414 327
rect 193 317 198 322
rect 409 317 414 322
rect 537 322 718 327
rect 801 322 1134 327
rect 1145 322 1214 327
rect 1329 322 1366 327
rect 1553 322 1678 327
rect 1745 322 2102 327
rect 2113 322 2158 327
rect 2193 322 2494 327
rect 2769 322 2870 327
rect 3137 322 3198 327
rect 3313 327 3318 332
rect 3313 322 3358 327
rect 537 317 542 322
rect 3137 317 3142 322
rect 105 312 150 317
rect 193 312 230 317
rect 273 312 302 317
rect 409 312 542 317
rect 601 312 742 317
rect 769 312 894 317
rect 1001 312 1334 317
rect 1353 312 1598 317
rect 1625 312 1942 317
rect 1993 312 2110 317
rect 2129 312 2390 317
rect 2409 312 2510 317
rect 2521 312 2582 317
rect 2705 312 2766 317
rect 2937 312 3142 317
rect 3169 312 3398 317
rect 273 307 278 312
rect 1329 307 1334 312
rect 2129 307 2134 312
rect 193 302 278 307
rect 313 302 342 307
rect 633 302 702 307
rect 761 302 918 307
rect 953 302 1110 307
rect 1329 302 1470 307
rect 1545 302 2134 307
rect 2385 307 2390 312
rect 2385 302 2758 307
rect 2873 302 2998 307
rect 3137 302 3254 307
rect 273 297 278 302
rect 1129 297 1254 302
rect 2169 297 2366 302
rect 2993 297 3078 302
rect 3137 297 3142 302
rect 273 292 302 297
rect 505 292 582 297
rect 745 292 878 297
rect 905 292 974 297
rect 1089 292 1134 297
rect 1249 292 1278 297
rect 1457 292 1606 297
rect 1673 292 1862 297
rect 1977 292 2118 297
rect 2145 292 2174 297
rect 2361 292 2566 297
rect 2665 292 2774 297
rect 2865 292 2974 297
rect 3073 292 3142 297
rect 297 287 390 292
rect 505 287 510 292
rect 385 277 390 287
rect 481 282 510 287
rect 577 287 582 292
rect 641 287 726 292
rect 577 282 646 287
rect 721 282 1174 287
rect 1185 282 1334 287
rect 1393 282 3054 287
rect 1185 277 1190 282
rect 153 272 366 277
rect 385 272 566 277
rect 657 272 1190 277
rect 1209 272 1374 277
rect 1465 272 2110 277
rect 2161 272 2478 277
rect 2785 272 2902 277
rect 153 267 158 272
rect 89 262 158 267
rect 361 267 366 272
rect 561 267 662 272
rect 2577 267 2694 272
rect 361 262 486 267
rect 681 262 782 267
rect 873 262 1230 267
rect 1489 262 1718 267
rect 1801 262 2062 267
rect 2073 262 2398 267
rect 2513 262 2582 267
rect 2689 262 2910 267
rect 1249 257 1358 262
rect 257 252 1110 257
rect 1161 252 1254 257
rect 1353 252 1598 257
rect 1641 252 2678 257
rect 2857 252 2886 257
rect 2673 247 2862 252
rect 169 242 374 247
rect 617 242 2126 247
rect 2345 242 2654 247
rect 2945 242 3038 247
rect 2121 237 2350 242
rect 2945 237 2950 242
rect 361 232 462 237
rect 521 232 1670 237
rect 1729 232 1854 237
rect 2369 232 2710 237
rect 2769 232 2950 237
rect 3033 237 3038 242
rect 3033 232 3286 237
rect 1873 227 2102 232
rect 2369 227 2374 232
rect 97 222 558 227
rect 673 222 822 227
rect 881 222 1654 227
rect 1665 222 1878 227
rect 2097 222 2374 227
rect 2385 222 2478 227
rect 2641 222 2670 227
rect 2473 217 2646 222
rect 177 212 214 217
rect 417 212 446 217
rect 441 207 446 212
rect 529 212 670 217
rect 529 207 534 212
rect 193 202 262 207
rect 441 202 534 207
rect 665 207 670 212
rect 769 212 990 217
rect 769 207 774 212
rect 665 202 774 207
rect 985 207 990 212
rect 1137 212 1406 217
rect 1137 207 1142 212
rect 1401 207 1406 212
rect 1497 212 1718 217
rect 1729 212 2078 217
rect 2105 212 2230 217
rect 2337 212 2454 217
rect 1497 207 1502 212
rect 985 202 1014 207
rect 1113 202 1142 207
rect 1201 202 1350 207
rect 1401 202 1502 207
rect 1713 207 1718 212
rect 2705 207 2710 232
rect 3033 222 3110 227
rect 3249 222 3318 227
rect 2745 212 2822 217
rect 2961 212 3078 217
rect 2961 207 2966 212
rect 3073 207 3078 212
rect 1713 202 2358 207
rect 2513 202 2598 207
rect 2705 202 2966 207
rect 2977 202 3054 207
rect 3073 202 3134 207
rect 3193 202 3270 207
rect 1009 197 1118 202
rect 1545 197 1694 202
rect 2513 197 2518 202
rect 185 192 342 197
rect 601 192 646 197
rect 793 192 870 197
rect 889 192 966 197
rect 1161 192 1382 197
rect 1521 192 1550 197
rect 1689 192 1934 197
rect 2041 192 2518 197
rect 2593 197 2598 202
rect 2593 192 2870 197
rect 3001 192 3118 197
rect 1953 187 2046 192
rect 553 182 814 187
rect 841 182 918 187
rect 985 182 1150 187
rect 1393 182 1582 187
rect 1593 182 1958 187
rect 2065 182 2366 187
rect 2377 182 2462 187
rect 2529 182 2582 187
rect 1145 177 1398 182
rect 2577 177 2582 182
rect 2769 182 2894 187
rect 2769 177 2774 182
rect 361 172 534 177
rect 553 172 622 177
rect 1657 172 1678 177
rect 1689 172 1830 177
rect 1945 172 2406 177
rect 2473 172 2558 177
rect 2577 172 2774 177
rect 2873 172 3206 177
rect 361 167 366 172
rect 281 162 366 167
rect 529 167 534 172
rect 641 167 846 172
rect 2401 167 2478 172
rect 529 162 646 167
rect 841 162 870 167
rect 1153 162 1278 167
rect 1297 162 1542 167
rect 1561 162 1830 167
rect 1881 162 1990 167
rect 2129 162 2382 167
rect 2793 162 2862 167
rect 1297 157 1302 162
rect 657 152 782 157
rect 833 152 902 157
rect 1065 152 1302 157
rect 1537 157 1542 162
rect 2009 157 2110 162
rect 2857 157 2862 162
rect 2921 162 2974 167
rect 2921 157 2926 162
rect 1537 152 2014 157
rect 2105 152 2502 157
rect 2577 152 2766 157
rect 2857 152 2926 157
rect 241 147 366 152
rect 657 147 662 152
rect 1329 147 1462 152
rect 2577 147 2582 152
rect 217 142 246 147
rect 361 142 662 147
rect 673 142 862 147
rect 921 142 1046 147
rect 921 137 926 142
rect 137 132 414 137
rect 561 132 694 137
rect 737 132 790 137
rect 809 132 926 137
rect 1041 137 1046 142
rect 1105 142 1334 147
rect 1457 142 1750 147
rect 1785 142 1926 147
rect 1953 142 2070 147
rect 2081 142 2582 147
rect 2761 147 2766 152
rect 2761 142 2790 147
rect 2945 142 3078 147
rect 3177 142 3302 147
rect 1105 137 1110 142
rect 1953 137 1958 142
rect 2601 137 2718 142
rect 1041 132 1110 137
rect 1129 132 1958 137
rect 1969 132 2254 137
rect 2297 132 2350 137
rect 2529 132 2606 137
rect 2713 132 2742 137
rect 2753 132 2814 137
rect 2833 132 2878 137
rect 409 127 566 132
rect 785 127 790 132
rect 2369 127 2510 132
rect 2833 127 2838 132
rect 2897 127 3030 132
rect 273 122 358 127
rect 593 122 702 127
rect 785 122 1494 127
rect 1505 122 1598 127
rect 1785 122 1814 127
rect 1825 122 2374 127
rect 2505 122 2838 127
rect 2857 122 2902 127
rect 3025 122 3102 127
rect 3281 122 3318 127
rect 1505 117 1510 122
rect 1593 117 1694 122
rect 1785 117 1790 122
rect 249 112 278 117
rect 273 107 278 112
rect 337 112 582 117
rect 337 107 342 112
rect 273 102 342 107
rect 577 107 582 112
rect 713 112 1510 117
rect 1537 112 1574 117
rect 1689 112 1790 117
rect 1809 117 1814 122
rect 1809 112 2118 117
rect 2137 112 2718 117
rect 713 107 718 112
rect 2113 107 2118 112
rect 2713 107 2718 112
rect 2801 112 3014 117
rect 2801 107 2806 112
rect 577 102 718 107
rect 745 102 966 107
rect 1121 102 1670 107
rect 1897 102 1982 107
rect 2113 102 2198 107
rect 2329 102 2694 107
rect 2713 102 2806 107
rect 2969 102 2998 107
rect 961 97 1126 102
rect 2001 97 2094 102
rect 2217 97 2310 102
rect 2993 97 2998 102
rect 3113 102 3310 107
rect 3113 97 3118 102
rect 361 92 390 97
rect 857 92 942 97
rect 1145 92 1430 97
rect 1521 92 2006 97
rect 2089 92 2222 97
rect 2305 92 2558 97
rect 2993 92 3118 97
rect 385 87 390 92
rect 761 87 862 92
rect 1425 87 1526 92
rect 2577 87 2702 92
rect 385 82 766 87
rect 1017 82 1166 87
rect 1337 82 1406 87
rect 1545 82 1638 87
rect 1905 82 2582 87
rect 2697 82 2942 87
rect 881 77 998 82
rect 1185 77 1318 82
rect 1681 77 1854 82
rect 785 72 886 77
rect 993 72 1190 77
rect 1313 72 1686 77
rect 1849 72 2686 77
rect 897 62 1406 67
rect 1513 62 1606 67
rect 1401 57 1518 62
rect 1601 57 1606 62
rect 1697 62 1838 67
rect 1953 62 2310 67
rect 2321 62 2414 67
rect 2513 62 2566 67
rect 2601 62 2822 67
rect 1697 57 1702 62
rect 1833 57 1958 62
rect 2513 57 2518 62
rect 777 52 1030 57
rect 1177 52 1382 57
rect 1025 47 1182 52
rect 1377 47 1382 52
rect 1537 52 1566 57
rect 1601 52 1702 57
rect 1977 52 2150 57
rect 2241 52 2518 57
rect 1537 47 1542 52
rect 1745 47 1814 52
rect 2705 47 2910 52
rect 849 42 1006 47
rect 1001 37 1006 42
rect 1201 42 1278 47
rect 1377 42 1542 47
rect 1721 42 1750 47
rect 1809 42 1926 47
rect 1985 42 2366 47
rect 2529 42 2710 47
rect 2905 42 2934 47
rect 1201 37 1206 42
rect 953 32 982 37
rect 1001 32 1206 37
rect 1225 32 1254 37
rect 977 17 982 32
rect 1225 17 1230 32
rect 1273 27 1278 42
rect 1721 37 1726 42
rect 2361 37 2534 42
rect 1577 32 1726 37
rect 1753 32 1798 37
rect 1577 27 1582 32
rect 1273 22 1582 27
rect 1793 27 1798 32
rect 2009 32 2190 37
rect 2313 32 2342 37
rect 2009 27 2014 32
rect 2337 27 2342 32
rect 2721 32 2798 37
rect 2721 27 2726 32
rect 1793 22 2014 27
rect 2033 22 2166 27
rect 2337 22 2726 27
rect 2793 27 2798 32
rect 2857 32 2886 37
rect 2857 27 2862 32
rect 2793 22 2862 27
rect 977 12 1230 17
rect 1745 12 1774 17
rect 1769 7 1774 12
rect 2201 12 2302 17
rect 2201 7 2206 12
rect 1769 2 2206 7
rect 2297 7 2302 12
rect 2745 12 2774 17
rect 2745 7 2750 12
rect 2297 2 2750 7
use AND2X2  AND2X2_0
timestamp 1711653199
transform 1 0 2880 0 -1 2170
box -8 -3 40 105
use AND2X2  AND2X2_1
timestamp 1711653199
transform 1 0 2712 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1711653199
transform 1 0 2592 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_3
timestamp 1711653199
transform 1 0 2704 0 1 2170
box -8 -3 40 105
use AND2X2  AND2X2_4
timestamp 1711653199
transform 1 0 288 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_5
timestamp 1711653199
transform 1 0 1160 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_6
timestamp 1711653199
transform 1 0 2576 0 -1 1170
box -8 -3 40 105
use AND2X2  AND2X2_7
timestamp 1711653199
transform 1 0 1880 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_8
timestamp 1711653199
transform 1 0 2096 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_9
timestamp 1711653199
transform 1 0 2032 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_10
timestamp 1711653199
transform 1 0 1856 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_11
timestamp 1711653199
transform 1 0 528 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_12
timestamp 1711653199
transform 1 0 192 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_13
timestamp 1711653199
transform 1 0 256 0 -1 1970
box -8 -3 40 105
use AND2X2  AND2X2_14
timestamp 1711653199
transform 1 0 104 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_15
timestamp 1711653199
transform 1 0 384 0 1 970
box -8 -3 40 105
use AND2X2  AND2X2_16
timestamp 1711653199
transform 1 0 656 0 -1 1570
box -8 -3 40 105
use AND2X2  AND2X2_17
timestamp 1711653199
transform 1 0 560 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_18
timestamp 1711653199
transform 1 0 544 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_19
timestamp 1711653199
transform 1 0 736 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_20
timestamp 1711653199
transform 1 0 904 0 1 1970
box -8 -3 40 105
use AND2X2  AND2X2_21
timestamp 1711653199
transform 1 0 680 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_22
timestamp 1711653199
transform 1 0 392 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_23
timestamp 1711653199
transform 1 0 368 0 -1 1970
box -8 -3 40 105
use AND2X2  AND2X2_24
timestamp 1711653199
transform 1 0 288 0 -1 370
box -8 -3 40 105
use AND2X2  AND2X2_25
timestamp 1711653199
transform 1 0 232 0 -1 2170
box -8 -3 40 105
use AND2X2  AND2X2_26
timestamp 1711653199
transform 1 0 1392 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_27
timestamp 1711653199
transform 1 0 944 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_28
timestamp 1711653199
transform 1 0 1160 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_29
timestamp 1711653199
transform 1 0 1200 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_30
timestamp 1711653199
transform 1 0 1136 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_31
timestamp 1711653199
transform 1 0 1152 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_32
timestamp 1711653199
transform 1 0 1080 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_33
timestamp 1711653199
transform 1 0 1952 0 -1 170
box -8 -3 40 105
use AND2X2  AND2X2_34
timestamp 1711653199
transform 1 0 2216 0 -1 770
box -8 -3 40 105
use AND2X2  AND2X2_35
timestamp 1711653199
transform 1 0 3280 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_36
timestamp 1711653199
transform 1 0 3240 0 1 1570
box -8 -3 40 105
use AND2X2  AND2X2_37
timestamp 1711653199
transform 1 0 3328 0 1 570
box -8 -3 40 105
use AND2X2  AND2X2_38
timestamp 1711653199
transform 1 0 3240 0 -1 1770
box -8 -3 40 105
use AND2X2  AND2X2_39
timestamp 1711653199
transform 1 0 2864 0 -1 370
box -8 -3 40 105
use AND2X2  AND2X2_40
timestamp 1711653199
transform 1 0 2768 0 1 1770
box -8 -3 40 105
use AND2X2  AND2X2_41
timestamp 1711653199
transform 1 0 2168 0 -1 2970
box -8 -3 40 105
use AND2X2  AND2X2_42
timestamp 1711653199
transform 1 0 832 0 -1 2970
box -8 -3 40 105
use AND2X2  AND2X2_43
timestamp 1711653199
transform 1 0 992 0 -1 2970
box -8 -3 40 105
use AND2X2  AND2X2_44
timestamp 1711653199
transform 1 0 1328 0 1 2970
box -8 -3 40 105
use AND2X2  AND2X2_45
timestamp 1711653199
transform 1 0 1512 0 -1 2970
box -8 -3 40 105
use AND2X2  AND2X2_46
timestamp 1711653199
transform 1 0 1248 0 -1 2970
box -8 -3 40 105
use AND2X2  AND2X2_47
timestamp 1711653199
transform 1 0 2776 0 -1 3170
box -8 -3 40 105
use AND2X2  AND2X2_48
timestamp 1711653199
transform 1 0 2464 0 1 2770
box -8 -3 40 105
use AND2X2  AND2X2_49
timestamp 1711653199
transform 1 0 2608 0 1 2770
box -8 -3 40 105
use AND2X2  AND2X2_50
timestamp 1711653199
transform 1 0 2912 0 1 2970
box -8 -3 40 105
use AND2X2  AND2X2_51
timestamp 1711653199
transform 1 0 2920 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_52
timestamp 1711653199
transform 1 0 3088 0 1 2170
box -8 -3 40 105
use AND2X2  AND2X2_53
timestamp 1711653199
transform 1 0 3288 0 -1 2170
box -8 -3 40 105
use AND2X2  AND2X2_54
timestamp 1711653199
transform 1 0 2840 0 -1 2370
box -8 -3 40 105
use AND2X2  AND2X2_55
timestamp 1711653199
transform 1 0 2784 0 1 2370
box -8 -3 40 105
use AND2X2  AND2X2_56
timestamp 1711653199
transform 1 0 2816 0 1 2770
box -8 -3 40 105
use AND2X2  AND2X2_57
timestamp 1711653199
transform 1 0 3024 0 -1 2770
box -8 -3 40 105
use AOI21X1  AOI21X1_0
timestamp 1711653199
transform 1 0 3024 0 1 2570
box -7 -3 39 105
use AOI21X1  AOI21X1_1
timestamp 1711653199
transform 1 0 2784 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_2
timestamp 1711653199
transform 1 0 2288 0 1 970
box -7 -3 39 105
use AOI21X1  AOI21X1_3
timestamp 1711653199
transform 1 0 2328 0 1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_4
timestamp 1711653199
transform 1 0 1752 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_5
timestamp 1711653199
transform 1 0 3048 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_6
timestamp 1711653199
transform 1 0 1024 0 1 1570
box -7 -3 39 105
use AOI21X1  AOI21X1_7
timestamp 1711653199
transform 1 0 2216 0 -1 1370
box -7 -3 39 105
use AOI21X1  AOI21X1_8
timestamp 1711653199
transform 1 0 2320 0 -1 370
box -7 -3 39 105
use AOI21X1  AOI21X1_9
timestamp 1711653199
transform 1 0 2464 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_10
timestamp 1711653199
transform 1 0 96 0 -1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_11
timestamp 1711653199
transform 1 0 2208 0 1 1170
box -7 -3 39 105
use AOI21X1  AOI21X1_12
timestamp 1711653199
transform 1 0 2088 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_13
timestamp 1711653199
transform 1 0 664 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_14
timestamp 1711653199
transform 1 0 432 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_15
timestamp 1711653199
transform 1 0 224 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_16
timestamp 1711653199
transform 1 0 344 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_17
timestamp 1711653199
transform 1 0 848 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_18
timestamp 1711653199
transform 1 0 2160 0 1 170
box -7 -3 39 105
use AOI21X1  AOI21X1_19
timestamp 1711653199
transform 1 0 2192 0 1 570
box -7 -3 39 105
use AOI21X1  AOI21X1_20
timestamp 1711653199
transform 1 0 776 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_21
timestamp 1711653199
transform 1 0 520 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_22
timestamp 1711653199
transform 1 0 352 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_23
timestamp 1711653199
transform 1 0 1352 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_24
timestamp 1711653199
transform 1 0 1928 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_25
timestamp 1711653199
transform 1 0 1728 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_26
timestamp 1711653199
transform 1 0 1816 0 1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_27
timestamp 1711653199
transform 1 0 3128 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_28
timestamp 1711653199
transform 1 0 3136 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_29
timestamp 1711653199
transform 1 0 3096 0 -1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_30
timestamp 1711653199
transform 1 0 2688 0 1 770
box -7 -3 39 105
use AOI21X1  AOI21X1_31
timestamp 1711653199
transform 1 0 2664 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_32
timestamp 1711653199
transform 1 0 2608 0 -1 2170
box -7 -3 39 105
use AOI21X1  AOI21X1_33
timestamp 1711653199
transform 1 0 2904 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_34
timestamp 1711653199
transform 1 0 3000 0 1 1970
box -7 -3 39 105
use AOI21X1  AOI21X1_35
timestamp 1711653199
transform 1 0 2624 0 1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_36
timestamp 1711653199
transform 1 0 2336 0 1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_37
timestamp 1711653199
transform 1 0 2472 0 1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_38
timestamp 1711653199
transform 1 0 2280 0 1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_39
timestamp 1711653199
transform 1 0 1008 0 1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_40
timestamp 1711653199
transform 1 0 1072 0 -1 2970
box -7 -3 39 105
use AOI21X1  AOI21X1_41
timestamp 1711653199
transform 1 0 952 0 -1 2770
box -7 -3 39 105
use AOI21X1  AOI21X1_42
timestamp 1711653199
transform 1 0 912 0 -1 2770
box -7 -3 39 105
use AOI22X1  AOI22X1_0
timestamp 1711653199
transform 1 0 2392 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_1
timestamp 1711653199
transform 1 0 2264 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_2
timestamp 1711653199
transform 1 0 2144 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_3
timestamp 1711653199
transform 1 0 2056 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_4
timestamp 1711653199
transform 1 0 3280 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_5
timestamp 1711653199
transform 1 0 952 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_6
timestamp 1711653199
transform 1 0 1224 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_7
timestamp 1711653199
transform 1 0 280 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_8
timestamp 1711653199
transform 1 0 704 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_9
timestamp 1711653199
transform 1 0 328 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_10
timestamp 1711653199
transform 1 0 288 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_11
timestamp 1711653199
transform 1 0 624 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_12
timestamp 1711653199
transform 1 0 392 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1711653199
transform 1 0 280 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_14
timestamp 1711653199
transform 1 0 1016 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_15
timestamp 1711653199
transform 1 0 1232 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_16
timestamp 1711653199
transform 1 0 264 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_17
timestamp 1711653199
transform 1 0 3288 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_18
timestamp 1711653199
transform 1 0 2056 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_19
timestamp 1711653199
transform 1 0 2248 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_20
timestamp 1711653199
transform 1 0 2464 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_21
timestamp 1711653199
transform 1 0 2536 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_22
timestamp 1711653199
transform 1 0 1904 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_23
timestamp 1711653199
transform 1 0 3336 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_24
timestamp 1711653199
transform 1 0 856 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_25
timestamp 1711653199
transform 1 0 1224 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_26
timestamp 1711653199
transform 1 0 288 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_27
timestamp 1711653199
transform 1 0 752 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_28
timestamp 1711653199
transform 1 0 424 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_29
timestamp 1711653199
transform 1 0 184 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_30
timestamp 1711653199
transform 1 0 1824 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_31
timestamp 1711653199
transform 1 0 1992 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_32
timestamp 1711653199
transform 1 0 2168 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_33
timestamp 1711653199
transform 1 0 976 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_34
timestamp 1711653199
transform 1 0 1208 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_35
timestamp 1711653199
transform 1 0 1936 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_36
timestamp 1711653199
transform 1 0 1856 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_37
timestamp 1711653199
transform 1 0 288 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_38
timestamp 1711653199
transform 1 0 2224 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_39
timestamp 1711653199
transform 1 0 1632 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_40
timestamp 1711653199
transform 1 0 3104 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_41
timestamp 1711653199
transform 1 0 1152 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_42
timestamp 1711653199
transform 1 0 520 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_43
timestamp 1711653199
transform 1 0 1632 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_44
timestamp 1711653199
transform 1 0 616 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_45
timestamp 1711653199
transform 1 0 384 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_46
timestamp 1711653199
transform 1 0 288 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1711653199
transform 1 0 936 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_48
timestamp 1711653199
transform 1 0 1152 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_49
timestamp 1711653199
transform 1 0 344 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_50
timestamp 1711653199
transform 1 0 3168 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_51
timestamp 1711653199
transform 1 0 2440 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_52
timestamp 1711653199
transform 1 0 1080 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_53
timestamp 1711653199
transform 1 0 520 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_54
timestamp 1711653199
transform 1 0 120 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_55
timestamp 1711653199
transform 1 0 2264 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_56
timestamp 1711653199
transform 1 0 1592 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_57
timestamp 1711653199
transform 1 0 3200 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_58
timestamp 1711653199
transform 1 0 912 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_59
timestamp 1711653199
transform 1 0 1216 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_60
timestamp 1711653199
transform 1 0 2008 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_61
timestamp 1711653199
transform 1 0 1856 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_62
timestamp 1711653199
transform 1 0 832 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_63
timestamp 1711653199
transform 1 0 1496 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_64
timestamp 1711653199
transform 1 0 1800 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_65
timestamp 1711653199
transform 1 0 176 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_66
timestamp 1711653199
transform 1 0 1648 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_67
timestamp 1711653199
transform 1 0 3104 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_68
timestamp 1711653199
transform 1 0 1264 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_69
timestamp 1711653199
transform 1 0 880 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_70
timestamp 1711653199
transform 1 0 864 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_71
timestamp 1711653199
transform 1 0 1392 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_72
timestamp 1711653199
transform 1 0 2424 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_73
timestamp 1711653199
transform 1 0 2512 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_74
timestamp 1711653199
transform 1 0 2024 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_75
timestamp 1711653199
transform 1 0 88 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_76
timestamp 1711653199
transform 1 0 2832 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_77
timestamp 1711653199
transform 1 0 3192 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_78
timestamp 1711653199
transform 1 0 1432 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_79
timestamp 1711653199
transform 1 0 472 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_80
timestamp 1711653199
transform 1 0 2080 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_81
timestamp 1711653199
transform 1 0 2408 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_82
timestamp 1711653199
transform 1 0 2248 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_83
timestamp 1711653199
transform 1 0 2480 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_84
timestamp 1711653199
transform 1 0 2304 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_85
timestamp 1711653199
transform 1 0 2568 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_86
timestamp 1711653199
transform 1 0 1992 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_87
timestamp 1711653199
transform 1 0 1896 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_88
timestamp 1711653199
transform 1 0 2384 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_89
timestamp 1711653199
transform 1 0 2312 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_90
timestamp 1711653199
transform 1 0 1960 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_91
timestamp 1711653199
transform 1 0 1848 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_92
timestamp 1711653199
transform 1 0 1880 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_93
timestamp 1711653199
transform 1 0 1656 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_94
timestamp 1711653199
transform 1 0 1616 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_95
timestamp 1711653199
transform 1 0 1736 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_96
timestamp 1711653199
transform 1 0 1616 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_97
timestamp 1711653199
transform 1 0 1528 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_98
timestamp 1711653199
transform 1 0 2120 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_99
timestamp 1711653199
transform 1 0 1920 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_100
timestamp 1711653199
transform 1 0 1896 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_101
timestamp 1711653199
transform 1 0 632 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_102
timestamp 1711653199
transform 1 0 616 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_103
timestamp 1711653199
transform 1 0 600 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_104
timestamp 1711653199
transform 1 0 600 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_105
timestamp 1711653199
transform 1 0 208 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_106
timestamp 1711653199
transform 1 0 208 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_107
timestamp 1711653199
transform 1 0 192 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_108
timestamp 1711653199
transform 1 0 224 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_109
timestamp 1711653199
transform 1 0 136 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_110
timestamp 1711653199
transform 1 0 160 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_111
timestamp 1711653199
transform 1 0 136 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_112
timestamp 1711653199
transform 1 0 88 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_113
timestamp 1711653199
transform 1 0 144 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_114
timestamp 1711653199
transform 1 0 336 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_115
timestamp 1711653199
transform 1 0 216 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_116
timestamp 1711653199
transform 1 0 192 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_117
timestamp 1711653199
transform 1 0 448 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_118
timestamp 1711653199
transform 1 0 600 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_119
timestamp 1711653199
transform 1 0 400 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_120
timestamp 1711653199
transform 1 0 496 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_121
timestamp 1711653199
transform 1 0 552 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_122
timestamp 1711653199
transform 1 0 680 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_123
timestamp 1711653199
transform 1 0 2248 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_124
timestamp 1711653199
transform 1 0 1696 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_125
timestamp 1711653199
transform 1 0 1800 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_126
timestamp 1711653199
transform 1 0 768 0 1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_127
timestamp 1711653199
transform 1 0 776 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_128
timestamp 1711653199
transform 1 0 760 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_129
timestamp 1711653199
transform 1 0 744 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_130
timestamp 1711653199
transform 1 0 856 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_131
timestamp 1711653199
transform 1 0 352 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_132
timestamp 1711653199
transform 1 0 344 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_133
timestamp 1711653199
transform 1 0 432 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_134
timestamp 1711653199
transform 1 0 336 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_135
timestamp 1711653199
transform 1 0 200 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_136
timestamp 1711653199
transform 1 0 288 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_137
timestamp 1711653199
transform 1 0 176 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_138
timestamp 1711653199
transform 1 0 96 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_139
timestamp 1711653199
transform 1 0 1344 0 1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_140
timestamp 1711653199
transform 1 0 1392 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_141
timestamp 1711653199
transform 1 0 1320 0 -1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_142
timestamp 1711653199
transform 1 0 1328 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_143
timestamp 1711653199
transform 1 0 1080 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_144
timestamp 1711653199
transform 1 0 936 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_145
timestamp 1711653199
transform 1 0 1280 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_146
timestamp 1711653199
transform 1 0 1224 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_147
timestamp 1711653199
transform 1 0 1032 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_148
timestamp 1711653199
transform 1 0 992 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_149
timestamp 1711653199
transform 1 0 2472 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_150
timestamp 1711653199
transform 1 0 2528 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_151
timestamp 1711653199
transform 1 0 1960 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_152
timestamp 1711653199
transform 1 0 1576 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_153
timestamp 1711653199
transform 1 0 3128 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_154
timestamp 1711653199
transform 1 0 2960 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_155
timestamp 1711653199
transform 1 0 3088 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_156
timestamp 1711653199
transform 1 0 3264 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_157
timestamp 1711653199
transform 1 0 3256 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_158
timestamp 1711653199
transform 1 0 3192 0 -1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_159
timestamp 1711653199
transform 1 0 3280 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_160
timestamp 1711653199
transform 1 0 3240 0 -1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_161
timestamp 1711653199
transform 1 0 3224 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_162
timestamp 1711653199
transform 1 0 3168 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_163
timestamp 1711653199
transform 1 0 3296 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_164
timestamp 1711653199
transform 1 0 2608 0 1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_165
timestamp 1711653199
transform 1 0 2672 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_166
timestamp 1711653199
transform 1 0 2728 0 1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_167
timestamp 1711653199
transform 1 0 2680 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_168
timestamp 1711653199
transform 1 0 2696 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_169
timestamp 1711653199
transform 1 0 2600 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_170
timestamp 1711653199
transform 1 0 2808 0 1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_171
timestamp 1711653199
transform 1 0 2544 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_172
timestamp 1711653199
transform 1 0 2560 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_173
timestamp 1711653199
transform 1 0 2880 0 -1 1170
box -8 -3 46 105
use AOI22X1  AOI22X1_174
timestamp 1711653199
transform 1 0 2776 0 1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_175
timestamp 1711653199
transform 1 0 2776 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_176
timestamp 1711653199
transform 1 0 2928 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_177
timestamp 1711653199
transform 1 0 3032 0 -1 1970
box -8 -3 46 105
use AOI22X1  AOI22X1_178
timestamp 1711653199
transform 1 0 2952 0 -1 1770
box -8 -3 46 105
use AOI22X1  AOI22X1_179
timestamp 1711653199
transform 1 0 2736 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_180
timestamp 1711653199
transform 1 0 2744 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_181
timestamp 1711653199
transform 1 0 2880 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_182
timestamp 1711653199
transform 1 0 3080 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_183
timestamp 1711653199
transform 1 0 3144 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_184
timestamp 1711653199
transform 1 0 3296 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_185
timestamp 1711653199
transform 1 0 2520 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_186
timestamp 1711653199
transform 1 0 2088 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_187
timestamp 1711653199
transform 1 0 2464 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_188
timestamp 1711653199
transform 1 0 2344 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_189
timestamp 1711653199
transform 1 0 2024 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_190
timestamp 1711653199
transform 1 0 840 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_191
timestamp 1711653199
transform 1 0 776 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_192
timestamp 1711653199
transform 1 0 680 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_193
timestamp 1711653199
transform 1 0 720 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_194
timestamp 1711653199
transform 1 0 1000 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_195
timestamp 1711653199
transform 1 0 784 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_196
timestamp 1711653199
transform 1 0 824 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_197
timestamp 1711653199
transform 1 0 920 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_198
timestamp 1711653199
transform 1 0 3200 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_199
timestamp 1711653199
transform 1 0 1576 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_200
timestamp 1711653199
transform 1 0 1856 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_201
timestamp 1711653199
transform 1 0 1896 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_202
timestamp 1711653199
transform 1 0 2544 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_203
timestamp 1711653199
transform 1 0 2640 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_204
timestamp 1711653199
transform 1 0 2312 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_205
timestamp 1711653199
transform 1 0 2112 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_206
timestamp 1711653199
transform 1 0 2112 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_207
timestamp 1711653199
transform 1 0 2072 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_208
timestamp 1711653199
transform 1 0 2152 0 1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_209
timestamp 1711653199
transform 1 0 1880 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_210
timestamp 1711653199
transform 1 0 1600 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_211
timestamp 1711653199
transform 1 0 1272 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_212
timestamp 1711653199
transform 1 0 1184 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_213
timestamp 1711653199
transform 1 0 1120 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_214
timestamp 1711653199
transform 1 0 1080 0 1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_215
timestamp 1711653199
transform 1 0 328 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_216
timestamp 1711653199
transform 1 0 240 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_217
timestamp 1711653199
transform 1 0 200 0 -1 2570
box -8 -3 46 105
use AOI22X1  AOI22X1_218
timestamp 1711653199
transform 1 0 112 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_219
timestamp 1711653199
transform 1 0 2360 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_220
timestamp 1711653199
transform 1 0 464 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_221
timestamp 1711653199
transform 1 0 400 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_222
timestamp 1711653199
transform 1 0 536 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_223
timestamp 1711653199
transform 1 0 856 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_224
timestamp 1711653199
transform 1 0 920 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_225
timestamp 1711653199
transform 1 0 600 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_226
timestamp 1711653199
transform 1 0 792 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_227
timestamp 1711653199
transform 1 0 1336 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_228
timestamp 1711653199
transform 1 0 1400 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_229
timestamp 1711653199
transform 1 0 1624 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_230
timestamp 1711653199
transform 1 0 1960 0 -1 2770
box -8 -3 46 105
use BUFX2  BUFX2_0
timestamp 1711653199
transform 1 0 1784 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1711653199
transform 1 0 1760 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_2
timestamp 1711653199
transform 1 0 2504 0 1 970
box -5 -3 28 105
use BUFX2  BUFX2_3
timestamp 1711653199
transform 1 0 3168 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_4
timestamp 1711653199
transform 1 0 3048 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_5
timestamp 1711653199
transform 1 0 2976 0 -1 1570
box -5 -3 28 105
use BUFX2  BUFX2_6
timestamp 1711653199
transform 1 0 2424 0 -1 1770
box -5 -3 28 105
use BUFX2  BUFX2_7
timestamp 1711653199
transform 1 0 2968 0 1 1770
box -5 -3 28 105
use BUFX2  BUFX2_8
timestamp 1711653199
transform 1 0 2608 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_9
timestamp 1711653199
transform 1 0 2584 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_10
timestamp 1711653199
transform 1 0 3168 0 -1 1970
box -5 -3 28 105
use BUFX2  BUFX2_11
timestamp 1711653199
transform 1 0 2776 0 1 2970
box -5 -3 28 105
use BUFX2  BUFX2_12
timestamp 1711653199
transform 1 0 2752 0 -1 2970
box -5 -3 28 105
use BUFX2  BUFX2_13
timestamp 1711653199
transform 1 0 1880 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_14
timestamp 1711653199
transform 1 0 1832 0 1 2770
box -5 -3 28 105
use BUFX2  BUFX2_15
timestamp 1711653199
transform 1 0 1808 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_16
timestamp 1711653199
transform 1 0 1456 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_17
timestamp 1711653199
transform 1 0 1224 0 1 2370
box -5 -3 28 105
use BUFX2  BUFX2_18
timestamp 1711653199
transform 1 0 1448 0 1 2370
box -5 -3 28 105
use BUFX2  BUFX2_19
timestamp 1711653199
transform 1 0 2960 0 1 2370
box -5 -3 28 105
use BUFX2  BUFX2_20
timestamp 1711653199
transform 1 0 1832 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_21
timestamp 1711653199
transform 1 0 3120 0 -1 970
box -5 -3 28 105
use BUFX2  BUFX2_22
timestamp 1711653199
transform 1 0 2952 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_23
timestamp 1711653199
transform 1 0 2664 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_24
timestamp 1711653199
transform 1 0 1920 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_25
timestamp 1711653199
transform 1 0 2032 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_26
timestamp 1711653199
transform 1 0 1736 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_27
timestamp 1711653199
transform 1 0 2128 0 -1 2770
box -5 -3 28 105
use BUFX2  BUFX2_28
timestamp 1711653199
transform 1 0 1664 0 1 2770
box -5 -3 28 105
use BUFX2  BUFX2_29
timestamp 1711653199
transform 1 0 2056 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_30
timestamp 1711653199
transform 1 0 2704 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_31
timestamp 1711653199
transform 1 0 2928 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_32
timestamp 1711653199
transform 1 0 3096 0 1 1570
box -5 -3 28 105
use BUFX2  BUFX2_33
timestamp 1711653199
transform 1 0 2776 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_34
timestamp 1711653199
transform 1 0 2408 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_35
timestamp 1711653199
transform 1 0 2384 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_36
timestamp 1711653199
transform 1 0 2184 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_37
timestamp 1711653199
transform 1 0 2608 0 -1 570
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1711653199
transform 1 0 3208 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1711653199
transform 1 0 3304 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1711653199
transform 1 0 2968 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1711653199
transform 1 0 3256 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1711653199
transform 1 0 2584 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1711653199
transform 1 0 2632 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1711653199
transform 1 0 2800 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1711653199
transform 1 0 2992 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1711653199
transform 1 0 2992 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1711653199
transform 1 0 2552 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1711653199
transform 1 0 2488 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1711653199
transform 1 0 2440 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1711653199
transform 1 0 2456 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1711653199
transform 1 0 2600 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1711653199
transform 1 0 2864 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1711653199
transform 1 0 2832 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1711653199
transform 1 0 2856 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1711653199
transform 1 0 3152 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1711653199
transform 1 0 3056 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1711653199
transform 1 0 2968 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1711653199
transform 1 0 3184 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1711653199
transform 1 0 2128 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1711653199
transform 1 0 2024 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1711653199
transform 1 0 1920 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1711653199
transform 1 0 1776 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1711653199
transform 1 0 1504 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1711653199
transform 1 0 1344 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1711653199
transform 1 0 1144 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1711653199
transform 1 0 1032 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1711653199
transform 1 0 296 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1711653199
transform 1 0 184 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1711653199
transform 1 0 80 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1711653199
transform 1 0 80 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1711653199
transform 1 0 448 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1711653199
transform 1 0 400 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1711653199
transform 1 0 512 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1711653199
transform 1 0 800 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1711653199
transform 1 0 832 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1711653199
transform 1 0 568 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1711653199
transform 1 0 680 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1711653199
transform 1 0 1400 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1711653199
transform 1 0 1352 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1711653199
transform 1 0 1616 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1711653199
transform 1 0 1504 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1711653199
transform 1 0 2184 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1711653199
transform 1 0 2024 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1711653199
transform 1 0 2544 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1711653199
transform 1 0 2544 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1711653199
transform 1 0 2432 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1711653199
transform 1 0 2176 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1711653199
transform 1 0 2288 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1711653199
transform 1 0 2328 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1711653199
transform 1 0 2224 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1711653199
transform 1 0 1712 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1711653199
transform 1 0 1872 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1711653199
transform 1 0 1704 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1711653199
transform 1 0 1488 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1711653199
transform 1 0 1256 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1711653199
transform 1 0 776 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1711653199
transform 1 0 552 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1711653199
transform 1 0 264 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1711653199
transform 1 0 408 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1711653199
transform 1 0 80 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1711653199
transform 1 0 80 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1711653199
transform 1 0 296 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1711653199
transform 1 0 160 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1711653199
transform 1 0 304 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1711653199
transform 1 0 304 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1711653199
transform 1 0 456 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_69
timestamp 1711653199
transform 1 0 568 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1711653199
transform 1 0 1144 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1711653199
transform 1 0 864 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1711653199
transform 1 0 1008 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1711653199
transform 1 0 1280 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1711653199
transform 1 0 1384 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1711653199
transform 1 0 1648 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1711653199
transform 1 0 1520 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1711653199
transform 1 0 1752 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1711653199
transform 1 0 1880 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1711653199
transform 1 0 2432 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_80
timestamp 1711653199
transform 1 0 2512 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1711653199
transform 1 0 2208 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1711653199
transform 1 0 2080 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_83
timestamp 1711653199
transform 1 0 2480 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_84
timestamp 1711653199
transform 1 0 2328 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1711653199
transform 1 0 1984 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1711653199
transform 1 0 2704 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1711653199
transform 1 0 1952 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1711653199
transform 1 0 1848 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_89
timestamp 1711653199
transform 1 0 1768 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1711653199
transform 1 0 1496 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1711653199
transform 1 0 968 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1711653199
transform 1 0 720 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1711653199
transform 1 0 328 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1711653199
transform 1 0 408 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_95
timestamp 1711653199
transform 1 0 192 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1711653199
transform 1 0 80 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1711653199
transform 1 0 80 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1711653199
transform 1 0 80 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1711653199
transform 1 0 264 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_100
timestamp 1711653199
transform 1 0 368 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_101
timestamp 1711653199
transform 1 0 416 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1711653199
transform 1 0 680 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1711653199
transform 1 0 992 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1711653199
transform 1 0 568 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_105
timestamp 1711653199
transform 1 0 808 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1711653199
transform 1 0 1288 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_107
timestamp 1711653199
transform 1 0 1456 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_108
timestamp 1711653199
transform 1 0 1696 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1711653199
transform 1 0 1560 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1711653199
transform 1 0 1800 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1711653199
transform 1 0 1912 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1711653199
transform 1 0 2496 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1711653199
transform 1 0 2704 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1711653199
transform 1 0 2264 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1711653199
transform 1 0 2064 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_116
timestamp 1711653199
transform 1 0 2160 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_117
timestamp 1711653199
transform 1 0 2360 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_118
timestamp 1711653199
transform 1 0 1960 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1711653199
transform 1 0 2792 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_120
timestamp 1711653199
transform 1 0 2888 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1711653199
transform 1 0 2816 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_122
timestamp 1711653199
transform 1 0 2808 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_123
timestamp 1711653199
transform 1 0 2888 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_124
timestamp 1711653199
transform 1 0 3304 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_125
timestamp 1711653199
transform 1 0 3192 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_126
timestamp 1711653199
transform 1 0 3296 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_127
timestamp 1711653199
transform 1 0 2960 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_128
timestamp 1711653199
transform 1 0 3080 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_129
timestamp 1711653199
transform 1 0 3304 0 -1 2970
box -8 -3 104 105
use FILL  FILL_0
timestamp 1711653199
transform 1 0 3392 0 1 3170
box -8 -3 16 105
use FILL  FILL_1
timestamp 1711653199
transform 1 0 3288 0 1 3170
box -8 -3 16 105
use FILL  FILL_2
timestamp 1711653199
transform 1 0 3184 0 1 3170
box -8 -3 16 105
use FILL  FILL_3
timestamp 1711653199
transform 1 0 3176 0 1 3170
box -8 -3 16 105
use FILL  FILL_4
timestamp 1711653199
transform 1 0 3072 0 1 3170
box -8 -3 16 105
use FILL  FILL_5
timestamp 1711653199
transform 1 0 3064 0 1 3170
box -8 -3 16 105
use FILL  FILL_6
timestamp 1711653199
transform 1 0 3056 0 1 3170
box -8 -3 16 105
use FILL  FILL_7
timestamp 1711653199
transform 1 0 2952 0 1 3170
box -8 -3 16 105
use FILL  FILL_8
timestamp 1711653199
transform 1 0 2912 0 1 3170
box -8 -3 16 105
use FILL  FILL_9
timestamp 1711653199
transform 1 0 2808 0 1 3170
box -8 -3 16 105
use FILL  FILL_10
timestamp 1711653199
transform 1 0 2800 0 1 3170
box -8 -3 16 105
use FILL  FILL_11
timestamp 1711653199
transform 1 0 2696 0 1 3170
box -8 -3 16 105
use FILL  FILL_12
timestamp 1711653199
transform 1 0 2688 0 1 3170
box -8 -3 16 105
use FILL  FILL_13
timestamp 1711653199
transform 1 0 2584 0 1 3170
box -8 -3 16 105
use FILL  FILL_14
timestamp 1711653199
transform 1 0 2576 0 1 3170
box -8 -3 16 105
use FILL  FILL_15
timestamp 1711653199
transform 1 0 2456 0 1 3170
box -8 -3 16 105
use FILL  FILL_16
timestamp 1711653199
transform 1 0 2448 0 1 3170
box -8 -3 16 105
use FILL  FILL_17
timestamp 1711653199
transform 1 0 2440 0 1 3170
box -8 -3 16 105
use FILL  FILL_18
timestamp 1711653199
transform 1 0 2320 0 1 3170
box -8 -3 16 105
use FILL  FILL_19
timestamp 1711653199
transform 1 0 2200 0 1 3170
box -8 -3 16 105
use FILL  FILL_20
timestamp 1711653199
transform 1 0 2192 0 1 3170
box -8 -3 16 105
use FILL  FILL_21
timestamp 1711653199
transform 1 0 1976 0 1 3170
box -8 -3 16 105
use FILL  FILL_22
timestamp 1711653199
transform 1 0 1872 0 1 3170
box -8 -3 16 105
use FILL  FILL_23
timestamp 1711653199
transform 1 0 1864 0 1 3170
box -8 -3 16 105
use FILL  FILL_24
timestamp 1711653199
transform 1 0 1744 0 1 3170
box -8 -3 16 105
use FILL  FILL_25
timestamp 1711653199
transform 1 0 1640 0 1 3170
box -8 -3 16 105
use FILL  FILL_26
timestamp 1711653199
transform 1 0 1632 0 1 3170
box -8 -3 16 105
use FILL  FILL_27
timestamp 1711653199
transform 1 0 1512 0 1 3170
box -8 -3 16 105
use FILL  FILL_28
timestamp 1711653199
transform 1 0 1504 0 1 3170
box -8 -3 16 105
use FILL  FILL_29
timestamp 1711653199
transform 1 0 1496 0 1 3170
box -8 -3 16 105
use FILL  FILL_30
timestamp 1711653199
transform 1 0 1376 0 1 3170
box -8 -3 16 105
use FILL  FILL_31
timestamp 1711653199
transform 1 0 1256 0 1 3170
box -8 -3 16 105
use FILL  FILL_32
timestamp 1711653199
transform 1 0 1248 0 1 3170
box -8 -3 16 105
use FILL  FILL_33
timestamp 1711653199
transform 1 0 1240 0 1 3170
box -8 -3 16 105
use FILL  FILL_34
timestamp 1711653199
transform 1 0 1136 0 1 3170
box -8 -3 16 105
use FILL  FILL_35
timestamp 1711653199
transform 1 0 1112 0 1 3170
box -8 -3 16 105
use FILL  FILL_36
timestamp 1711653199
transform 1 0 1104 0 1 3170
box -8 -3 16 105
use FILL  FILL_37
timestamp 1711653199
transform 1 0 1000 0 1 3170
box -8 -3 16 105
use FILL  FILL_38
timestamp 1711653199
transform 1 0 976 0 1 3170
box -8 -3 16 105
use FILL  FILL_39
timestamp 1711653199
transform 1 0 968 0 1 3170
box -8 -3 16 105
use FILL  FILL_40
timestamp 1711653199
transform 1 0 960 0 1 3170
box -8 -3 16 105
use FILL  FILL_41
timestamp 1711653199
transform 1 0 856 0 1 3170
box -8 -3 16 105
use FILL  FILL_42
timestamp 1711653199
transform 1 0 848 0 1 3170
box -8 -3 16 105
use FILL  FILL_43
timestamp 1711653199
transform 1 0 840 0 1 3170
box -8 -3 16 105
use FILL  FILL_44
timestamp 1711653199
transform 1 0 832 0 1 3170
box -8 -3 16 105
use FILL  FILL_45
timestamp 1711653199
transform 1 0 808 0 1 3170
box -8 -3 16 105
use FILL  FILL_46
timestamp 1711653199
transform 1 0 800 0 1 3170
box -8 -3 16 105
use FILL  FILL_47
timestamp 1711653199
transform 1 0 792 0 1 3170
box -8 -3 16 105
use FILL  FILL_48
timestamp 1711653199
transform 1 0 784 0 1 3170
box -8 -3 16 105
use FILL  FILL_49
timestamp 1711653199
transform 1 0 752 0 1 3170
box -8 -3 16 105
use FILL  FILL_50
timestamp 1711653199
transform 1 0 744 0 1 3170
box -8 -3 16 105
use FILL  FILL_51
timestamp 1711653199
transform 1 0 688 0 1 3170
box -8 -3 16 105
use FILL  FILL_52
timestamp 1711653199
transform 1 0 680 0 1 3170
box -8 -3 16 105
use FILL  FILL_53
timestamp 1711653199
transform 1 0 672 0 1 3170
box -8 -3 16 105
use FILL  FILL_54
timestamp 1711653199
transform 1 0 664 0 1 3170
box -8 -3 16 105
use FILL  FILL_55
timestamp 1711653199
transform 1 0 560 0 1 3170
box -8 -3 16 105
use FILL  FILL_56
timestamp 1711653199
transform 1 0 552 0 1 3170
box -8 -3 16 105
use FILL  FILL_57
timestamp 1711653199
transform 1 0 448 0 1 3170
box -8 -3 16 105
use FILL  FILL_58
timestamp 1711653199
transform 1 0 424 0 1 3170
box -8 -3 16 105
use FILL  FILL_59
timestamp 1711653199
transform 1 0 416 0 1 3170
box -8 -3 16 105
use FILL  FILL_60
timestamp 1711653199
transform 1 0 408 0 1 3170
box -8 -3 16 105
use FILL  FILL_61
timestamp 1711653199
transform 1 0 400 0 1 3170
box -8 -3 16 105
use FILL  FILL_62
timestamp 1711653199
transform 1 0 296 0 1 3170
box -8 -3 16 105
use FILL  FILL_63
timestamp 1711653199
transform 1 0 288 0 1 3170
box -8 -3 16 105
use FILL  FILL_64
timestamp 1711653199
transform 1 0 264 0 1 3170
box -8 -3 16 105
use FILL  FILL_65
timestamp 1711653199
transform 1 0 256 0 1 3170
box -8 -3 16 105
use FILL  FILL_66
timestamp 1711653199
transform 1 0 152 0 1 3170
box -8 -3 16 105
use FILL  FILL_67
timestamp 1711653199
transform 1 0 144 0 1 3170
box -8 -3 16 105
use FILL  FILL_68
timestamp 1711653199
transform 1 0 136 0 1 3170
box -8 -3 16 105
use FILL  FILL_69
timestamp 1711653199
transform 1 0 128 0 1 3170
box -8 -3 16 105
use FILL  FILL_70
timestamp 1711653199
transform 1 0 120 0 1 3170
box -8 -3 16 105
use FILL  FILL_71
timestamp 1711653199
transform 1 0 112 0 1 3170
box -8 -3 16 105
use FILL  FILL_72
timestamp 1711653199
transform 1 0 104 0 1 3170
box -8 -3 16 105
use FILL  FILL_73
timestamp 1711653199
transform 1 0 96 0 1 3170
box -8 -3 16 105
use FILL  FILL_74
timestamp 1711653199
transform 1 0 88 0 1 3170
box -8 -3 16 105
use FILL  FILL_75
timestamp 1711653199
transform 1 0 80 0 1 3170
box -8 -3 16 105
use FILL  FILL_76
timestamp 1711653199
transform 1 0 72 0 1 3170
box -8 -3 16 105
use FILL  FILL_77
timestamp 1711653199
transform 1 0 3392 0 -1 3170
box -8 -3 16 105
use FILL  FILL_78
timestamp 1711653199
transform 1 0 3384 0 -1 3170
box -8 -3 16 105
use FILL  FILL_79
timestamp 1711653199
transform 1 0 3376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_80
timestamp 1711653199
transform 1 0 3368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_81
timestamp 1711653199
transform 1 0 3360 0 -1 3170
box -8 -3 16 105
use FILL  FILL_82
timestamp 1711653199
transform 1 0 3320 0 -1 3170
box -8 -3 16 105
use FILL  FILL_83
timestamp 1711653199
transform 1 0 3312 0 -1 3170
box -8 -3 16 105
use FILL  FILL_84
timestamp 1711653199
transform 1 0 3256 0 -1 3170
box -8 -3 16 105
use FILL  FILL_85
timestamp 1711653199
transform 1 0 3248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_86
timestamp 1711653199
transform 1 0 3240 0 -1 3170
box -8 -3 16 105
use FILL  FILL_87
timestamp 1711653199
transform 1 0 3232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_88
timestamp 1711653199
transform 1 0 3176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_89
timestamp 1711653199
transform 1 0 3168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_90
timestamp 1711653199
transform 1 0 3136 0 -1 3170
box -8 -3 16 105
use FILL  FILL_91
timestamp 1711653199
transform 1 0 3104 0 -1 3170
box -8 -3 16 105
use FILL  FILL_92
timestamp 1711653199
transform 1 0 3096 0 -1 3170
box -8 -3 16 105
use FILL  FILL_93
timestamp 1711653199
transform 1 0 3088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_94
timestamp 1711653199
transform 1 0 3032 0 -1 3170
box -8 -3 16 105
use FILL  FILL_95
timestamp 1711653199
transform 1 0 3024 0 -1 3170
box -8 -3 16 105
use FILL  FILL_96
timestamp 1711653199
transform 1 0 3000 0 -1 3170
box -8 -3 16 105
use FILL  FILL_97
timestamp 1711653199
transform 1 0 2992 0 -1 3170
box -8 -3 16 105
use FILL  FILL_98
timestamp 1711653199
transform 1 0 2984 0 -1 3170
box -8 -3 16 105
use FILL  FILL_99
timestamp 1711653199
transform 1 0 2880 0 -1 3170
box -8 -3 16 105
use FILL  FILL_100
timestamp 1711653199
transform 1 0 2872 0 -1 3170
box -8 -3 16 105
use FILL  FILL_101
timestamp 1711653199
transform 1 0 2864 0 -1 3170
box -8 -3 16 105
use FILL  FILL_102
timestamp 1711653199
transform 1 0 2832 0 -1 3170
box -8 -3 16 105
use FILL  FILL_103
timestamp 1711653199
transform 1 0 2824 0 -1 3170
box -8 -3 16 105
use FILL  FILL_104
timestamp 1711653199
transform 1 0 2768 0 -1 3170
box -8 -3 16 105
use FILL  FILL_105
timestamp 1711653199
transform 1 0 2760 0 -1 3170
box -8 -3 16 105
use FILL  FILL_106
timestamp 1711653199
transform 1 0 2696 0 -1 3170
box -8 -3 16 105
use FILL  FILL_107
timestamp 1711653199
transform 1 0 2688 0 -1 3170
box -8 -3 16 105
use FILL  FILL_108
timestamp 1711653199
transform 1 0 2632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_109
timestamp 1711653199
transform 1 0 2560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_110
timestamp 1711653199
transform 1 0 2552 0 -1 3170
box -8 -3 16 105
use FILL  FILL_111
timestamp 1711653199
transform 1 0 2544 0 -1 3170
box -8 -3 16 105
use FILL  FILL_112
timestamp 1711653199
transform 1 0 2456 0 -1 3170
box -8 -3 16 105
use FILL  FILL_113
timestamp 1711653199
transform 1 0 2448 0 -1 3170
box -8 -3 16 105
use FILL  FILL_114
timestamp 1711653199
transform 1 0 2440 0 -1 3170
box -8 -3 16 105
use FILL  FILL_115
timestamp 1711653199
transform 1 0 2432 0 -1 3170
box -8 -3 16 105
use FILL  FILL_116
timestamp 1711653199
transform 1 0 2352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_117
timestamp 1711653199
transform 1 0 2344 0 -1 3170
box -8 -3 16 105
use FILL  FILL_118
timestamp 1711653199
transform 1 0 2336 0 -1 3170
box -8 -3 16 105
use FILL  FILL_119
timestamp 1711653199
transform 1 0 2328 0 -1 3170
box -8 -3 16 105
use FILL  FILL_120
timestamp 1711653199
transform 1 0 2272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_121
timestamp 1711653199
transform 1 0 2248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_122
timestamp 1711653199
transform 1 0 2200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_123
timestamp 1711653199
transform 1 0 2192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_124
timestamp 1711653199
transform 1 0 2152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_125
timestamp 1711653199
transform 1 0 2120 0 -1 3170
box -8 -3 16 105
use FILL  FILL_126
timestamp 1711653199
transform 1 0 2080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_127
timestamp 1711653199
transform 1 0 2072 0 -1 3170
box -8 -3 16 105
use FILL  FILL_128
timestamp 1711653199
transform 1 0 2064 0 -1 3170
box -8 -3 16 105
use FILL  FILL_129
timestamp 1711653199
transform 1 0 2008 0 -1 3170
box -8 -3 16 105
use FILL  FILL_130
timestamp 1711653199
transform 1 0 2000 0 -1 3170
box -8 -3 16 105
use FILL  FILL_131
timestamp 1711653199
transform 1 0 1992 0 -1 3170
box -8 -3 16 105
use FILL  FILL_132
timestamp 1711653199
transform 1 0 1904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_133
timestamp 1711653199
transform 1 0 1896 0 -1 3170
box -8 -3 16 105
use FILL  FILL_134
timestamp 1711653199
transform 1 0 1888 0 -1 3170
box -8 -3 16 105
use FILL  FILL_135
timestamp 1711653199
transform 1 0 1880 0 -1 3170
box -8 -3 16 105
use FILL  FILL_136
timestamp 1711653199
transform 1 0 1848 0 -1 3170
box -8 -3 16 105
use FILL  FILL_137
timestamp 1711653199
transform 1 0 1776 0 -1 3170
box -8 -3 16 105
use FILL  FILL_138
timestamp 1711653199
transform 1 0 1768 0 -1 3170
box -8 -3 16 105
use FILL  FILL_139
timestamp 1711653199
transform 1 0 1760 0 -1 3170
box -8 -3 16 105
use FILL  FILL_140
timestamp 1711653199
transform 1 0 1752 0 -1 3170
box -8 -3 16 105
use FILL  FILL_141
timestamp 1711653199
transform 1 0 1672 0 -1 3170
box -8 -3 16 105
use FILL  FILL_142
timestamp 1711653199
transform 1 0 1664 0 -1 3170
box -8 -3 16 105
use FILL  FILL_143
timestamp 1711653199
transform 1 0 1656 0 -1 3170
box -8 -3 16 105
use FILL  FILL_144
timestamp 1711653199
transform 1 0 1648 0 -1 3170
box -8 -3 16 105
use FILL  FILL_145
timestamp 1711653199
transform 1 0 1640 0 -1 3170
box -8 -3 16 105
use FILL  FILL_146
timestamp 1711653199
transform 1 0 1576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_147
timestamp 1711653199
transform 1 0 1568 0 -1 3170
box -8 -3 16 105
use FILL  FILL_148
timestamp 1711653199
transform 1 0 1528 0 -1 3170
box -8 -3 16 105
use FILL  FILL_149
timestamp 1711653199
transform 1 0 1520 0 -1 3170
box -8 -3 16 105
use FILL  FILL_150
timestamp 1711653199
transform 1 0 1456 0 -1 3170
box -8 -3 16 105
use FILL  FILL_151
timestamp 1711653199
transform 1 0 1448 0 -1 3170
box -8 -3 16 105
use FILL  FILL_152
timestamp 1711653199
transform 1 0 1440 0 -1 3170
box -8 -3 16 105
use FILL  FILL_153
timestamp 1711653199
transform 1 0 1384 0 -1 3170
box -8 -3 16 105
use FILL  FILL_154
timestamp 1711653199
transform 1 0 1376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_155
timestamp 1711653199
transform 1 0 1336 0 -1 3170
box -8 -3 16 105
use FILL  FILL_156
timestamp 1711653199
transform 1 0 1272 0 -1 3170
box -8 -3 16 105
use FILL  FILL_157
timestamp 1711653199
transform 1 0 1264 0 -1 3170
box -8 -3 16 105
use FILL  FILL_158
timestamp 1711653199
transform 1 0 1232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_159
timestamp 1711653199
transform 1 0 1224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_160
timestamp 1711653199
transform 1 0 1152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_161
timestamp 1711653199
transform 1 0 1144 0 -1 3170
box -8 -3 16 105
use FILL  FILL_162
timestamp 1711653199
transform 1 0 1136 0 -1 3170
box -8 -3 16 105
use FILL  FILL_163
timestamp 1711653199
transform 1 0 1104 0 -1 3170
box -8 -3 16 105
use FILL  FILL_164
timestamp 1711653199
transform 1 0 1032 0 -1 3170
box -8 -3 16 105
use FILL  FILL_165
timestamp 1711653199
transform 1 0 1024 0 -1 3170
box -8 -3 16 105
use FILL  FILL_166
timestamp 1711653199
transform 1 0 1016 0 -1 3170
box -8 -3 16 105
use FILL  FILL_167
timestamp 1711653199
transform 1 0 1008 0 -1 3170
box -8 -3 16 105
use FILL  FILL_168
timestamp 1711653199
transform 1 0 912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_169
timestamp 1711653199
transform 1 0 904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_170
timestamp 1711653199
transform 1 0 800 0 -1 3170
box -8 -3 16 105
use FILL  FILL_171
timestamp 1711653199
transform 1 0 672 0 -1 3170
box -8 -3 16 105
use FILL  FILL_172
timestamp 1711653199
transform 1 0 664 0 -1 3170
box -8 -3 16 105
use FILL  FILL_173
timestamp 1711653199
transform 1 0 560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_174
timestamp 1711653199
transform 1 0 552 0 -1 3170
box -8 -3 16 105
use FILL  FILL_175
timestamp 1711653199
transform 1 0 544 0 -1 3170
box -8 -3 16 105
use FILL  FILL_176
timestamp 1711653199
transform 1 0 480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_177
timestamp 1711653199
transform 1 0 472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_178
timestamp 1711653199
transform 1 0 416 0 -1 3170
box -8 -3 16 105
use FILL  FILL_179
timestamp 1711653199
transform 1 0 408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_180
timestamp 1711653199
transform 1 0 400 0 -1 3170
box -8 -3 16 105
use FILL  FILL_181
timestamp 1711653199
transform 1 0 296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_182
timestamp 1711653199
transform 1 0 288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_183
timestamp 1711653199
transform 1 0 280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_184
timestamp 1711653199
transform 1 0 240 0 -1 3170
box -8 -3 16 105
use FILL  FILL_185
timestamp 1711653199
transform 1 0 232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_186
timestamp 1711653199
transform 1 0 176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_187
timestamp 1711653199
transform 1 0 168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_188
timestamp 1711653199
transform 1 0 160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_189
timestamp 1711653199
transform 1 0 152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_190
timestamp 1711653199
transform 1 0 144 0 -1 3170
box -8 -3 16 105
use FILL  FILL_191
timestamp 1711653199
transform 1 0 136 0 -1 3170
box -8 -3 16 105
use FILL  FILL_192
timestamp 1711653199
transform 1 0 128 0 -1 3170
box -8 -3 16 105
use FILL  FILL_193
timestamp 1711653199
transform 1 0 120 0 -1 3170
box -8 -3 16 105
use FILL  FILL_194
timestamp 1711653199
transform 1 0 112 0 -1 3170
box -8 -3 16 105
use FILL  FILL_195
timestamp 1711653199
transform 1 0 104 0 -1 3170
box -8 -3 16 105
use FILL  FILL_196
timestamp 1711653199
transform 1 0 96 0 -1 3170
box -8 -3 16 105
use FILL  FILL_197
timestamp 1711653199
transform 1 0 88 0 -1 3170
box -8 -3 16 105
use FILL  FILL_198
timestamp 1711653199
transform 1 0 80 0 -1 3170
box -8 -3 16 105
use FILL  FILL_199
timestamp 1711653199
transform 1 0 72 0 -1 3170
box -8 -3 16 105
use FILL  FILL_200
timestamp 1711653199
transform 1 0 3296 0 1 2970
box -8 -3 16 105
use FILL  FILL_201
timestamp 1711653199
transform 1 0 3288 0 1 2970
box -8 -3 16 105
use FILL  FILL_202
timestamp 1711653199
transform 1 0 3176 0 1 2970
box -8 -3 16 105
use FILL  FILL_203
timestamp 1711653199
transform 1 0 3168 0 1 2970
box -8 -3 16 105
use FILL  FILL_204
timestamp 1711653199
transform 1 0 3160 0 1 2970
box -8 -3 16 105
use FILL  FILL_205
timestamp 1711653199
transform 1 0 3152 0 1 2970
box -8 -3 16 105
use FILL  FILL_206
timestamp 1711653199
transform 1 0 3056 0 1 2970
box -8 -3 16 105
use FILL  FILL_207
timestamp 1711653199
transform 1 0 3048 0 1 2970
box -8 -3 16 105
use FILL  FILL_208
timestamp 1711653199
transform 1 0 3040 0 1 2970
box -8 -3 16 105
use FILL  FILL_209
timestamp 1711653199
transform 1 0 2968 0 1 2970
box -8 -3 16 105
use FILL  FILL_210
timestamp 1711653199
transform 1 0 2944 0 1 2970
box -8 -3 16 105
use FILL  FILL_211
timestamp 1711653199
transform 1 0 2904 0 1 2970
box -8 -3 16 105
use FILL  FILL_212
timestamp 1711653199
transform 1 0 2800 0 1 2970
box -8 -3 16 105
use FILL  FILL_213
timestamp 1711653199
transform 1 0 2696 0 1 2970
box -8 -3 16 105
use FILL  FILL_214
timestamp 1711653199
transform 1 0 2688 0 1 2970
box -8 -3 16 105
use FILL  FILL_215
timestamp 1711653199
transform 1 0 2680 0 1 2970
box -8 -3 16 105
use FILL  FILL_216
timestamp 1711653199
transform 1 0 2600 0 1 2970
box -8 -3 16 105
use FILL  FILL_217
timestamp 1711653199
transform 1 0 2592 0 1 2970
box -8 -3 16 105
use FILL  FILL_218
timestamp 1711653199
transform 1 0 2584 0 1 2970
box -8 -3 16 105
use FILL  FILL_219
timestamp 1711653199
transform 1 0 2576 0 1 2970
box -8 -3 16 105
use FILL  FILL_220
timestamp 1711653199
transform 1 0 2512 0 1 2970
box -8 -3 16 105
use FILL  FILL_221
timestamp 1711653199
transform 1 0 2504 0 1 2970
box -8 -3 16 105
use FILL  FILL_222
timestamp 1711653199
transform 1 0 2432 0 1 2970
box -8 -3 16 105
use FILL  FILL_223
timestamp 1711653199
transform 1 0 2424 0 1 2970
box -8 -3 16 105
use FILL  FILL_224
timestamp 1711653199
transform 1 0 2416 0 1 2970
box -8 -3 16 105
use FILL  FILL_225
timestamp 1711653199
transform 1 0 2392 0 1 2970
box -8 -3 16 105
use FILL  FILL_226
timestamp 1711653199
transform 1 0 2328 0 1 2970
box -8 -3 16 105
use FILL  FILL_227
timestamp 1711653199
transform 1 0 2320 0 1 2970
box -8 -3 16 105
use FILL  FILL_228
timestamp 1711653199
transform 1 0 2312 0 1 2970
box -8 -3 16 105
use FILL  FILL_229
timestamp 1711653199
transform 1 0 2256 0 1 2970
box -8 -3 16 105
use FILL  FILL_230
timestamp 1711653199
transform 1 0 2208 0 1 2970
box -8 -3 16 105
use FILL  FILL_231
timestamp 1711653199
transform 1 0 2200 0 1 2970
box -8 -3 16 105
use FILL  FILL_232
timestamp 1711653199
transform 1 0 2160 0 1 2970
box -8 -3 16 105
use FILL  FILL_233
timestamp 1711653199
transform 1 0 2152 0 1 2970
box -8 -3 16 105
use FILL  FILL_234
timestamp 1711653199
transform 1 0 2144 0 1 2970
box -8 -3 16 105
use FILL  FILL_235
timestamp 1711653199
transform 1 0 2080 0 1 2970
box -8 -3 16 105
use FILL  FILL_236
timestamp 1711653199
transform 1 0 2016 0 1 2970
box -8 -3 16 105
use FILL  FILL_237
timestamp 1711653199
transform 1 0 2008 0 1 2970
box -8 -3 16 105
use FILL  FILL_238
timestamp 1711653199
transform 1 0 1904 0 1 2970
box -8 -3 16 105
use FILL  FILL_239
timestamp 1711653199
transform 1 0 1816 0 1 2970
box -8 -3 16 105
use FILL  FILL_240
timestamp 1711653199
transform 1 0 1808 0 1 2970
box -8 -3 16 105
use FILL  FILL_241
timestamp 1711653199
transform 1 0 1800 0 1 2970
box -8 -3 16 105
use FILL  FILL_242
timestamp 1711653199
transform 1 0 1728 0 1 2970
box -8 -3 16 105
use FILL  FILL_243
timestamp 1711653199
transform 1 0 1664 0 1 2970
box -8 -3 16 105
use FILL  FILL_244
timestamp 1711653199
transform 1 0 1656 0 1 2970
box -8 -3 16 105
use FILL  FILL_245
timestamp 1711653199
transform 1 0 1592 0 1 2970
box -8 -3 16 105
use FILL  FILL_246
timestamp 1711653199
transform 1 0 1584 0 1 2970
box -8 -3 16 105
use FILL  FILL_247
timestamp 1711653199
transform 1 0 1536 0 1 2970
box -8 -3 16 105
use FILL  FILL_248
timestamp 1711653199
transform 1 0 1472 0 1 2970
box -8 -3 16 105
use FILL  FILL_249
timestamp 1711653199
transform 1 0 1464 0 1 2970
box -8 -3 16 105
use FILL  FILL_250
timestamp 1711653199
transform 1 0 1456 0 1 2970
box -8 -3 16 105
use FILL  FILL_251
timestamp 1711653199
transform 1 0 1432 0 1 2970
box -8 -3 16 105
use FILL  FILL_252
timestamp 1711653199
transform 1 0 1360 0 1 2970
box -8 -3 16 105
use FILL  FILL_253
timestamp 1711653199
transform 1 0 1280 0 1 2970
box -8 -3 16 105
use FILL  FILL_254
timestamp 1711653199
transform 1 0 1272 0 1 2970
box -8 -3 16 105
use FILL  FILL_255
timestamp 1711653199
transform 1 0 1184 0 1 2970
box -8 -3 16 105
use FILL  FILL_256
timestamp 1711653199
transform 1 0 1176 0 1 2970
box -8 -3 16 105
use FILL  FILL_257
timestamp 1711653199
transform 1 0 1168 0 1 2970
box -8 -3 16 105
use FILL  FILL_258
timestamp 1711653199
transform 1 0 1088 0 1 2970
box -8 -3 16 105
use FILL  FILL_259
timestamp 1711653199
transform 1 0 1040 0 1 2970
box -8 -3 16 105
use FILL  FILL_260
timestamp 1711653199
transform 1 0 1000 0 1 2970
box -8 -3 16 105
use FILL  FILL_261
timestamp 1711653199
transform 1 0 952 0 1 2970
box -8 -3 16 105
use FILL  FILL_262
timestamp 1711653199
transform 1 0 912 0 1 2970
box -8 -3 16 105
use FILL  FILL_263
timestamp 1711653199
transform 1 0 904 0 1 2970
box -8 -3 16 105
use FILL  FILL_264
timestamp 1711653199
transform 1 0 896 0 1 2970
box -8 -3 16 105
use FILL  FILL_265
timestamp 1711653199
transform 1 0 832 0 1 2970
box -8 -3 16 105
use FILL  FILL_266
timestamp 1711653199
transform 1 0 768 0 1 2970
box -8 -3 16 105
use FILL  FILL_267
timestamp 1711653199
transform 1 0 760 0 1 2970
box -8 -3 16 105
use FILL  FILL_268
timestamp 1711653199
transform 1 0 672 0 1 2970
box -8 -3 16 105
use FILL  FILL_269
timestamp 1711653199
transform 1 0 664 0 1 2970
box -8 -3 16 105
use FILL  FILL_270
timestamp 1711653199
transform 1 0 600 0 1 2970
box -8 -3 16 105
use FILL  FILL_271
timestamp 1711653199
transform 1 0 592 0 1 2970
box -8 -3 16 105
use FILL  FILL_272
timestamp 1711653199
transform 1 0 520 0 1 2970
box -8 -3 16 105
use FILL  FILL_273
timestamp 1711653199
transform 1 0 512 0 1 2970
box -8 -3 16 105
use FILL  FILL_274
timestamp 1711653199
transform 1 0 408 0 1 2970
box -8 -3 16 105
use FILL  FILL_275
timestamp 1711653199
transform 1 0 376 0 1 2970
box -8 -3 16 105
use FILL  FILL_276
timestamp 1711653199
transform 1 0 368 0 1 2970
box -8 -3 16 105
use FILL  FILL_277
timestamp 1711653199
transform 1 0 360 0 1 2970
box -8 -3 16 105
use FILL  FILL_278
timestamp 1711653199
transform 1 0 280 0 1 2970
box -8 -3 16 105
use FILL  FILL_279
timestamp 1711653199
transform 1 0 272 0 1 2970
box -8 -3 16 105
use FILL  FILL_280
timestamp 1711653199
transform 1 0 264 0 1 2970
box -8 -3 16 105
use FILL  FILL_281
timestamp 1711653199
transform 1 0 232 0 1 2970
box -8 -3 16 105
use FILL  FILL_282
timestamp 1711653199
transform 1 0 184 0 1 2970
box -8 -3 16 105
use FILL  FILL_283
timestamp 1711653199
transform 1 0 176 0 1 2970
box -8 -3 16 105
use FILL  FILL_284
timestamp 1711653199
transform 1 0 72 0 1 2970
box -8 -3 16 105
use FILL  FILL_285
timestamp 1711653199
transform 1 0 3296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_286
timestamp 1711653199
transform 1 0 3288 0 -1 2970
box -8 -3 16 105
use FILL  FILL_287
timestamp 1711653199
transform 1 0 3192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_288
timestamp 1711653199
transform 1 0 3184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_289
timestamp 1711653199
transform 1 0 3176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_290
timestamp 1711653199
transform 1 0 3096 0 -1 2970
box -8 -3 16 105
use FILL  FILL_291
timestamp 1711653199
transform 1 0 3088 0 -1 2970
box -8 -3 16 105
use FILL  FILL_292
timestamp 1711653199
transform 1 0 2992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_293
timestamp 1711653199
transform 1 0 2984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_294
timestamp 1711653199
transform 1 0 2784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_295
timestamp 1711653199
transform 1 0 2776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_296
timestamp 1711653199
transform 1 0 2696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_297
timestamp 1711653199
transform 1 0 2688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_298
timestamp 1711653199
transform 1 0 2608 0 -1 2970
box -8 -3 16 105
use FILL  FILL_299
timestamp 1711653199
transform 1 0 2504 0 -1 2970
box -8 -3 16 105
use FILL  FILL_300
timestamp 1711653199
transform 1 0 2424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_301
timestamp 1711653199
transform 1 0 2416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_302
timestamp 1711653199
transform 1 0 2312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_303
timestamp 1711653199
transform 1 0 2304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_304
timestamp 1711653199
transform 1 0 2208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_305
timestamp 1711653199
transform 1 0 2200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_306
timestamp 1711653199
transform 1 0 2128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_307
timestamp 1711653199
transform 1 0 2088 0 -1 2970
box -8 -3 16 105
use FILL  FILL_308
timestamp 1711653199
transform 1 0 2016 0 -1 2970
box -8 -3 16 105
use FILL  FILL_309
timestamp 1711653199
transform 1 0 2008 0 -1 2970
box -8 -3 16 105
use FILL  FILL_310
timestamp 1711653199
transform 1 0 2000 0 -1 2970
box -8 -3 16 105
use FILL  FILL_311
timestamp 1711653199
transform 1 0 1992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_312
timestamp 1711653199
transform 1 0 1912 0 -1 2970
box -8 -3 16 105
use FILL  FILL_313
timestamp 1711653199
transform 1 0 1792 0 -1 2970
box -8 -3 16 105
use FILL  FILL_314
timestamp 1711653199
transform 1 0 1688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_315
timestamp 1711653199
transform 1 0 1552 0 -1 2970
box -8 -3 16 105
use FILL  FILL_316
timestamp 1711653199
transform 1 0 1544 0 -1 2970
box -8 -3 16 105
use FILL  FILL_317
timestamp 1711653199
transform 1 0 1472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_318
timestamp 1711653199
transform 1 0 1464 0 -1 2970
box -8 -3 16 105
use FILL  FILL_319
timestamp 1711653199
transform 1 0 1424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_320
timestamp 1711653199
transform 1 0 1360 0 -1 2970
box -8 -3 16 105
use FILL  FILL_321
timestamp 1711653199
transform 1 0 1352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_322
timestamp 1711653199
transform 1 0 1344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_323
timestamp 1711653199
transform 1 0 1280 0 -1 2970
box -8 -3 16 105
use FILL  FILL_324
timestamp 1711653199
transform 1 0 1224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_325
timestamp 1711653199
transform 1 0 1216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_326
timestamp 1711653199
transform 1 0 1152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_327
timestamp 1711653199
transform 1 0 1144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_328
timestamp 1711653199
transform 1 0 1064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_329
timestamp 1711653199
transform 1 0 1056 0 -1 2970
box -8 -3 16 105
use FILL  FILL_330
timestamp 1711653199
transform 1 0 1032 0 -1 2970
box -8 -3 16 105
use FILL  FILL_331
timestamp 1711653199
transform 1 0 1024 0 -1 2970
box -8 -3 16 105
use FILL  FILL_332
timestamp 1711653199
transform 1 0 928 0 -1 2970
box -8 -3 16 105
use FILL  FILL_333
timestamp 1711653199
transform 1 0 920 0 -1 2970
box -8 -3 16 105
use FILL  FILL_334
timestamp 1711653199
transform 1 0 912 0 -1 2970
box -8 -3 16 105
use FILL  FILL_335
timestamp 1711653199
transform 1 0 792 0 -1 2970
box -8 -3 16 105
use FILL  FILL_336
timestamp 1711653199
transform 1 0 784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_337
timestamp 1711653199
transform 1 0 776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_338
timestamp 1711653199
transform 1 0 696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_339
timestamp 1711653199
transform 1 0 672 0 -1 2970
box -8 -3 16 105
use FILL  FILL_340
timestamp 1711653199
transform 1 0 664 0 -1 2970
box -8 -3 16 105
use FILL  FILL_341
timestamp 1711653199
transform 1 0 656 0 -1 2970
box -8 -3 16 105
use FILL  FILL_342
timestamp 1711653199
transform 1 0 592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_343
timestamp 1711653199
transform 1 0 584 0 -1 2970
box -8 -3 16 105
use FILL  FILL_344
timestamp 1711653199
transform 1 0 544 0 -1 2970
box -8 -3 16 105
use FILL  FILL_345
timestamp 1711653199
transform 1 0 536 0 -1 2970
box -8 -3 16 105
use FILL  FILL_346
timestamp 1711653199
transform 1 0 472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_347
timestamp 1711653199
transform 1 0 464 0 -1 2970
box -8 -3 16 105
use FILL  FILL_348
timestamp 1711653199
transform 1 0 360 0 -1 2970
box -8 -3 16 105
use FILL  FILL_349
timestamp 1711653199
transform 1 0 256 0 -1 2970
box -8 -3 16 105
use FILL  FILL_350
timestamp 1711653199
transform 1 0 248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_351
timestamp 1711653199
transform 1 0 184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_352
timestamp 1711653199
transform 1 0 176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_353
timestamp 1711653199
transform 1 0 72 0 -1 2970
box -8 -3 16 105
use FILL  FILL_354
timestamp 1711653199
transform 1 0 3392 0 1 2770
box -8 -3 16 105
use FILL  FILL_355
timestamp 1711653199
transform 1 0 3336 0 1 2770
box -8 -3 16 105
use FILL  FILL_356
timestamp 1711653199
transform 1 0 3264 0 1 2770
box -8 -3 16 105
use FILL  FILL_357
timestamp 1711653199
transform 1 0 3256 0 1 2770
box -8 -3 16 105
use FILL  FILL_358
timestamp 1711653199
transform 1 0 3248 0 1 2770
box -8 -3 16 105
use FILL  FILL_359
timestamp 1711653199
transform 1 0 3240 0 1 2770
box -8 -3 16 105
use FILL  FILL_360
timestamp 1711653199
transform 1 0 3168 0 1 2770
box -8 -3 16 105
use FILL  FILL_361
timestamp 1711653199
transform 1 0 3160 0 1 2770
box -8 -3 16 105
use FILL  FILL_362
timestamp 1711653199
transform 1 0 3152 0 1 2770
box -8 -3 16 105
use FILL  FILL_363
timestamp 1711653199
transform 1 0 3144 0 1 2770
box -8 -3 16 105
use FILL  FILL_364
timestamp 1711653199
transform 1 0 3136 0 1 2770
box -8 -3 16 105
use FILL  FILL_365
timestamp 1711653199
transform 1 0 3080 0 1 2770
box -8 -3 16 105
use FILL  FILL_366
timestamp 1711653199
transform 1 0 3072 0 1 2770
box -8 -3 16 105
use FILL  FILL_367
timestamp 1711653199
transform 1 0 3040 0 1 2770
box -8 -3 16 105
use FILL  FILL_368
timestamp 1711653199
transform 1 0 3032 0 1 2770
box -8 -3 16 105
use FILL  FILL_369
timestamp 1711653199
transform 1 0 3024 0 1 2770
box -8 -3 16 105
use FILL  FILL_370
timestamp 1711653199
transform 1 0 2968 0 1 2770
box -8 -3 16 105
use FILL  FILL_371
timestamp 1711653199
transform 1 0 2960 0 1 2770
box -8 -3 16 105
use FILL  FILL_372
timestamp 1711653199
transform 1 0 2952 0 1 2770
box -8 -3 16 105
use FILL  FILL_373
timestamp 1711653199
transform 1 0 2848 0 1 2770
box -8 -3 16 105
use FILL  FILL_374
timestamp 1711653199
transform 1 0 2808 0 1 2770
box -8 -3 16 105
use FILL  FILL_375
timestamp 1711653199
transform 1 0 2800 0 1 2770
box -8 -3 16 105
use FILL  FILL_376
timestamp 1711653199
transform 1 0 2696 0 1 2770
box -8 -3 16 105
use FILL  FILL_377
timestamp 1711653199
transform 1 0 2688 0 1 2770
box -8 -3 16 105
use FILL  FILL_378
timestamp 1711653199
transform 1 0 2680 0 1 2770
box -8 -3 16 105
use FILL  FILL_379
timestamp 1711653199
transform 1 0 2600 0 1 2770
box -8 -3 16 105
use FILL  FILL_380
timestamp 1711653199
transform 1 0 2592 0 1 2770
box -8 -3 16 105
use FILL  FILL_381
timestamp 1711653199
transform 1 0 2456 0 1 2770
box -8 -3 16 105
use FILL  FILL_382
timestamp 1711653199
transform 1 0 2256 0 1 2770
box -8 -3 16 105
use FILL  FILL_383
timestamp 1711653199
transform 1 0 2056 0 1 2770
box -8 -3 16 105
use FILL  FILL_384
timestamp 1711653199
transform 1 0 1952 0 1 2770
box -8 -3 16 105
use FILL  FILL_385
timestamp 1711653199
transform 1 0 1944 0 1 2770
box -8 -3 16 105
use FILL  FILL_386
timestamp 1711653199
transform 1 0 1936 0 1 2770
box -8 -3 16 105
use FILL  FILL_387
timestamp 1711653199
transform 1 0 1824 0 1 2770
box -8 -3 16 105
use FILL  FILL_388
timestamp 1711653199
transform 1 0 1816 0 1 2770
box -8 -3 16 105
use FILL  FILL_389
timestamp 1711653199
transform 1 0 1808 0 1 2770
box -8 -3 16 105
use FILL  FILL_390
timestamp 1711653199
transform 1 0 1704 0 1 2770
box -8 -3 16 105
use FILL  FILL_391
timestamp 1711653199
transform 1 0 1696 0 1 2770
box -8 -3 16 105
use FILL  FILL_392
timestamp 1711653199
transform 1 0 1688 0 1 2770
box -8 -3 16 105
use FILL  FILL_393
timestamp 1711653199
transform 1 0 1616 0 1 2770
box -8 -3 16 105
use FILL  FILL_394
timestamp 1711653199
transform 1 0 1568 0 1 2770
box -8 -3 16 105
use FILL  FILL_395
timestamp 1711653199
transform 1 0 1560 0 1 2770
box -8 -3 16 105
use FILL  FILL_396
timestamp 1711653199
transform 1 0 1552 0 1 2770
box -8 -3 16 105
use FILL  FILL_397
timestamp 1711653199
transform 1 0 1448 0 1 2770
box -8 -3 16 105
use FILL  FILL_398
timestamp 1711653199
transform 1 0 1440 0 1 2770
box -8 -3 16 105
use FILL  FILL_399
timestamp 1711653199
transform 1 0 1392 0 1 2770
box -8 -3 16 105
use FILL  FILL_400
timestamp 1711653199
transform 1 0 1384 0 1 2770
box -8 -3 16 105
use FILL  FILL_401
timestamp 1711653199
transform 1 0 1280 0 1 2770
box -8 -3 16 105
use FILL  FILL_402
timestamp 1711653199
transform 1 0 1272 0 1 2770
box -8 -3 16 105
use FILL  FILL_403
timestamp 1711653199
transform 1 0 1264 0 1 2770
box -8 -3 16 105
use FILL  FILL_404
timestamp 1711653199
transform 1 0 1256 0 1 2770
box -8 -3 16 105
use FILL  FILL_405
timestamp 1711653199
transform 1 0 1224 0 1 2770
box -8 -3 16 105
use FILL  FILL_406
timestamp 1711653199
transform 1 0 1152 0 1 2770
box -8 -3 16 105
use FILL  FILL_407
timestamp 1711653199
transform 1 0 1144 0 1 2770
box -8 -3 16 105
use FILL  FILL_408
timestamp 1711653199
transform 1 0 1136 0 1 2770
box -8 -3 16 105
use FILL  FILL_409
timestamp 1711653199
transform 1 0 1128 0 1 2770
box -8 -3 16 105
use FILL  FILL_410
timestamp 1711653199
transform 1 0 1120 0 1 2770
box -8 -3 16 105
use FILL  FILL_411
timestamp 1711653199
transform 1 0 1096 0 1 2770
box -8 -3 16 105
use FILL  FILL_412
timestamp 1711653199
transform 1 0 1088 0 1 2770
box -8 -3 16 105
use FILL  FILL_413
timestamp 1711653199
transform 1 0 984 0 1 2770
box -8 -3 16 105
use FILL  FILL_414
timestamp 1711653199
transform 1 0 976 0 1 2770
box -8 -3 16 105
use FILL  FILL_415
timestamp 1711653199
transform 1 0 968 0 1 2770
box -8 -3 16 105
use FILL  FILL_416
timestamp 1711653199
transform 1 0 960 0 1 2770
box -8 -3 16 105
use FILL  FILL_417
timestamp 1711653199
transform 1 0 912 0 1 2770
box -8 -3 16 105
use FILL  FILL_418
timestamp 1711653199
transform 1 0 904 0 1 2770
box -8 -3 16 105
use FILL  FILL_419
timestamp 1711653199
transform 1 0 896 0 1 2770
box -8 -3 16 105
use FILL  FILL_420
timestamp 1711653199
transform 1 0 848 0 1 2770
box -8 -3 16 105
use FILL  FILL_421
timestamp 1711653199
transform 1 0 840 0 1 2770
box -8 -3 16 105
use FILL  FILL_422
timestamp 1711653199
transform 1 0 832 0 1 2770
box -8 -3 16 105
use FILL  FILL_423
timestamp 1711653199
transform 1 0 784 0 1 2770
box -8 -3 16 105
use FILL  FILL_424
timestamp 1711653199
transform 1 0 776 0 1 2770
box -8 -3 16 105
use FILL  FILL_425
timestamp 1711653199
transform 1 0 768 0 1 2770
box -8 -3 16 105
use FILL  FILL_426
timestamp 1711653199
transform 1 0 760 0 1 2770
box -8 -3 16 105
use FILL  FILL_427
timestamp 1711653199
transform 1 0 712 0 1 2770
box -8 -3 16 105
use FILL  FILL_428
timestamp 1711653199
transform 1 0 704 0 1 2770
box -8 -3 16 105
use FILL  FILL_429
timestamp 1711653199
transform 1 0 696 0 1 2770
box -8 -3 16 105
use FILL  FILL_430
timestamp 1711653199
transform 1 0 648 0 1 2770
box -8 -3 16 105
use FILL  FILL_431
timestamp 1711653199
transform 1 0 640 0 1 2770
box -8 -3 16 105
use FILL  FILL_432
timestamp 1711653199
transform 1 0 592 0 1 2770
box -8 -3 16 105
use FILL  FILL_433
timestamp 1711653199
transform 1 0 584 0 1 2770
box -8 -3 16 105
use FILL  FILL_434
timestamp 1711653199
transform 1 0 576 0 1 2770
box -8 -3 16 105
use FILL  FILL_435
timestamp 1711653199
transform 1 0 528 0 1 2770
box -8 -3 16 105
use FILL  FILL_436
timestamp 1711653199
transform 1 0 520 0 1 2770
box -8 -3 16 105
use FILL  FILL_437
timestamp 1711653199
transform 1 0 512 0 1 2770
box -8 -3 16 105
use FILL  FILL_438
timestamp 1711653199
transform 1 0 504 0 1 2770
box -8 -3 16 105
use FILL  FILL_439
timestamp 1711653199
transform 1 0 456 0 1 2770
box -8 -3 16 105
use FILL  FILL_440
timestamp 1711653199
transform 1 0 448 0 1 2770
box -8 -3 16 105
use FILL  FILL_441
timestamp 1711653199
transform 1 0 440 0 1 2770
box -8 -3 16 105
use FILL  FILL_442
timestamp 1711653199
transform 1 0 392 0 1 2770
box -8 -3 16 105
use FILL  FILL_443
timestamp 1711653199
transform 1 0 384 0 1 2770
box -8 -3 16 105
use FILL  FILL_444
timestamp 1711653199
transform 1 0 376 0 1 2770
box -8 -3 16 105
use FILL  FILL_445
timestamp 1711653199
transform 1 0 368 0 1 2770
box -8 -3 16 105
use FILL  FILL_446
timestamp 1711653199
transform 1 0 320 0 1 2770
box -8 -3 16 105
use FILL  FILL_447
timestamp 1711653199
transform 1 0 312 0 1 2770
box -8 -3 16 105
use FILL  FILL_448
timestamp 1711653199
transform 1 0 304 0 1 2770
box -8 -3 16 105
use FILL  FILL_449
timestamp 1711653199
transform 1 0 296 0 1 2770
box -8 -3 16 105
use FILL  FILL_450
timestamp 1711653199
transform 1 0 288 0 1 2770
box -8 -3 16 105
use FILL  FILL_451
timestamp 1711653199
transform 1 0 184 0 1 2770
box -8 -3 16 105
use FILL  FILL_452
timestamp 1711653199
transform 1 0 176 0 1 2770
box -8 -3 16 105
use FILL  FILL_453
timestamp 1711653199
transform 1 0 168 0 1 2770
box -8 -3 16 105
use FILL  FILL_454
timestamp 1711653199
transform 1 0 160 0 1 2770
box -8 -3 16 105
use FILL  FILL_455
timestamp 1711653199
transform 1 0 152 0 1 2770
box -8 -3 16 105
use FILL  FILL_456
timestamp 1711653199
transform 1 0 104 0 1 2770
box -8 -3 16 105
use FILL  FILL_457
timestamp 1711653199
transform 1 0 96 0 1 2770
box -8 -3 16 105
use FILL  FILL_458
timestamp 1711653199
transform 1 0 88 0 1 2770
box -8 -3 16 105
use FILL  FILL_459
timestamp 1711653199
transform 1 0 80 0 1 2770
box -8 -3 16 105
use FILL  FILL_460
timestamp 1711653199
transform 1 0 72 0 1 2770
box -8 -3 16 105
use FILL  FILL_461
timestamp 1711653199
transform 1 0 3392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_462
timestamp 1711653199
transform 1 0 3384 0 -1 2770
box -8 -3 16 105
use FILL  FILL_463
timestamp 1711653199
transform 1 0 3280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_464
timestamp 1711653199
transform 1 0 3016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_465
timestamp 1711653199
transform 1 0 2928 0 -1 2770
box -8 -3 16 105
use FILL  FILL_466
timestamp 1711653199
transform 1 0 2920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_467
timestamp 1711653199
transform 1 0 2888 0 -1 2770
box -8 -3 16 105
use FILL  FILL_468
timestamp 1711653199
transform 1 0 2800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_469
timestamp 1711653199
transform 1 0 2792 0 -1 2770
box -8 -3 16 105
use FILL  FILL_470
timestamp 1711653199
transform 1 0 2704 0 -1 2770
box -8 -3 16 105
use FILL  FILL_471
timestamp 1711653199
transform 1 0 2696 0 -1 2770
box -8 -3 16 105
use FILL  FILL_472
timestamp 1711653199
transform 1 0 2592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_473
timestamp 1711653199
transform 1 0 2584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_474
timestamp 1711653199
transform 1 0 2536 0 -1 2770
box -8 -3 16 105
use FILL  FILL_475
timestamp 1711653199
transform 1 0 2528 0 -1 2770
box -8 -3 16 105
use FILL  FILL_476
timestamp 1711653199
transform 1 0 2424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_477
timestamp 1711653199
transform 1 0 2416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_478
timestamp 1711653199
transform 1 0 2408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_479
timestamp 1711653199
transform 1 0 2400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_480
timestamp 1711653199
transform 1 0 2352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_481
timestamp 1711653199
transform 1 0 2304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_482
timestamp 1711653199
transform 1 0 2296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_483
timestamp 1711653199
transform 1 0 2288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_484
timestamp 1711653199
transform 1 0 2280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_485
timestamp 1711653199
transform 1 0 2176 0 -1 2770
box -8 -3 16 105
use FILL  FILL_486
timestamp 1711653199
transform 1 0 2168 0 -1 2770
box -8 -3 16 105
use FILL  FILL_487
timestamp 1711653199
transform 1 0 2120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_488
timestamp 1711653199
transform 1 0 2016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_489
timestamp 1711653199
transform 1 0 2008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_490
timestamp 1711653199
transform 1 0 2000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_491
timestamp 1711653199
transform 1 0 1952 0 -1 2770
box -8 -3 16 105
use FILL  FILL_492
timestamp 1711653199
transform 1 0 1944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_493
timestamp 1711653199
transform 1 0 1872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_494
timestamp 1711653199
transform 1 0 1864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_495
timestamp 1711653199
transform 1 0 1856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_496
timestamp 1711653199
transform 1 0 1728 0 -1 2770
box -8 -3 16 105
use FILL  FILL_497
timestamp 1711653199
transform 1 0 1720 0 -1 2770
box -8 -3 16 105
use FILL  FILL_498
timestamp 1711653199
transform 1 0 1712 0 -1 2770
box -8 -3 16 105
use FILL  FILL_499
timestamp 1711653199
transform 1 0 1608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_500
timestamp 1711653199
transform 1 0 1600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_501
timestamp 1711653199
transform 1 0 1496 0 -1 2770
box -8 -3 16 105
use FILL  FILL_502
timestamp 1711653199
transform 1 0 1392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_503
timestamp 1711653199
transform 1 0 1384 0 -1 2770
box -8 -3 16 105
use FILL  FILL_504
timestamp 1711653199
transform 1 0 1376 0 -1 2770
box -8 -3 16 105
use FILL  FILL_505
timestamp 1711653199
transform 1 0 1328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_506
timestamp 1711653199
transform 1 0 1320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_507
timestamp 1711653199
transform 1 0 1280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_508
timestamp 1711653199
transform 1 0 1272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_509
timestamp 1711653199
transform 1 0 1224 0 -1 2770
box -8 -3 16 105
use FILL  FILL_510
timestamp 1711653199
transform 1 0 1216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_511
timestamp 1711653199
transform 1 0 1152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_512
timestamp 1711653199
transform 1 0 1112 0 -1 2770
box -8 -3 16 105
use FILL  FILL_513
timestamp 1711653199
transform 1 0 1104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_514
timestamp 1711653199
transform 1 0 1096 0 -1 2770
box -8 -3 16 105
use FILL  FILL_515
timestamp 1711653199
transform 1 0 1024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_516
timestamp 1711653199
transform 1 0 1016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_517
timestamp 1711653199
transform 1 0 1008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_518
timestamp 1711653199
transform 1 0 1000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_519
timestamp 1711653199
transform 1 0 944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_520
timestamp 1711653199
transform 1 0 888 0 -1 2770
box -8 -3 16 105
use FILL  FILL_521
timestamp 1711653199
transform 1 0 880 0 -1 2770
box -8 -3 16 105
use FILL  FILL_522
timestamp 1711653199
transform 1 0 872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_523
timestamp 1711653199
transform 1 0 864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_524
timestamp 1711653199
transform 1 0 800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_525
timestamp 1711653199
transform 1 0 792 0 -1 2770
box -8 -3 16 105
use FILL  FILL_526
timestamp 1711653199
transform 1 0 728 0 -1 2770
box -8 -3 16 105
use FILL  FILL_527
timestamp 1711653199
transform 1 0 720 0 -1 2770
box -8 -3 16 105
use FILL  FILL_528
timestamp 1711653199
transform 1 0 712 0 -1 2770
box -8 -3 16 105
use FILL  FILL_529
timestamp 1711653199
transform 1 0 704 0 -1 2770
box -8 -3 16 105
use FILL  FILL_530
timestamp 1711653199
transform 1 0 696 0 -1 2770
box -8 -3 16 105
use FILL  FILL_531
timestamp 1711653199
transform 1 0 608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_532
timestamp 1711653199
transform 1 0 600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_533
timestamp 1711653199
transform 1 0 592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_534
timestamp 1711653199
transform 1 0 584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_535
timestamp 1711653199
transform 1 0 520 0 -1 2770
box -8 -3 16 105
use FILL  FILL_536
timestamp 1711653199
transform 1 0 488 0 -1 2770
box -8 -3 16 105
use FILL  FILL_537
timestamp 1711653199
transform 1 0 480 0 -1 2770
box -8 -3 16 105
use FILL  FILL_538
timestamp 1711653199
transform 1 0 472 0 -1 2770
box -8 -3 16 105
use FILL  FILL_539
timestamp 1711653199
transform 1 0 400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_540
timestamp 1711653199
transform 1 0 392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_541
timestamp 1711653199
transform 1 0 288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_542
timestamp 1711653199
transform 1 0 280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_543
timestamp 1711653199
transform 1 0 272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_544
timestamp 1711653199
transform 1 0 264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_545
timestamp 1711653199
transform 1 0 192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_546
timestamp 1711653199
transform 1 0 184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_547
timestamp 1711653199
transform 1 0 176 0 -1 2770
box -8 -3 16 105
use FILL  FILL_548
timestamp 1711653199
transform 1 0 72 0 -1 2770
box -8 -3 16 105
use FILL  FILL_549
timestamp 1711653199
transform 1 0 3392 0 1 2570
box -8 -3 16 105
use FILL  FILL_550
timestamp 1711653199
transform 1 0 3384 0 1 2570
box -8 -3 16 105
use FILL  FILL_551
timestamp 1711653199
transform 1 0 3336 0 1 2570
box -8 -3 16 105
use FILL  FILL_552
timestamp 1711653199
transform 1 0 3288 0 1 2570
box -8 -3 16 105
use FILL  FILL_553
timestamp 1711653199
transform 1 0 3280 0 1 2570
box -8 -3 16 105
use FILL  FILL_554
timestamp 1711653199
transform 1 0 3232 0 1 2570
box -8 -3 16 105
use FILL  FILL_555
timestamp 1711653199
transform 1 0 3224 0 1 2570
box -8 -3 16 105
use FILL  FILL_556
timestamp 1711653199
transform 1 0 3216 0 1 2570
box -8 -3 16 105
use FILL  FILL_557
timestamp 1711653199
transform 1 0 3208 0 1 2570
box -8 -3 16 105
use FILL  FILL_558
timestamp 1711653199
transform 1 0 3200 0 1 2570
box -8 -3 16 105
use FILL  FILL_559
timestamp 1711653199
transform 1 0 3136 0 1 2570
box -8 -3 16 105
use FILL  FILL_560
timestamp 1711653199
transform 1 0 3128 0 1 2570
box -8 -3 16 105
use FILL  FILL_561
timestamp 1711653199
transform 1 0 3120 0 1 2570
box -8 -3 16 105
use FILL  FILL_562
timestamp 1711653199
transform 1 0 3072 0 1 2570
box -8 -3 16 105
use FILL  FILL_563
timestamp 1711653199
transform 1 0 3016 0 1 2570
box -8 -3 16 105
use FILL  FILL_564
timestamp 1711653199
transform 1 0 3008 0 1 2570
box -8 -3 16 105
use FILL  FILL_565
timestamp 1711653199
transform 1 0 3000 0 1 2570
box -8 -3 16 105
use FILL  FILL_566
timestamp 1711653199
transform 1 0 2992 0 1 2570
box -8 -3 16 105
use FILL  FILL_567
timestamp 1711653199
transform 1 0 2928 0 1 2570
box -8 -3 16 105
use FILL  FILL_568
timestamp 1711653199
transform 1 0 2920 0 1 2570
box -8 -3 16 105
use FILL  FILL_569
timestamp 1711653199
transform 1 0 2856 0 1 2570
box -8 -3 16 105
use FILL  FILL_570
timestamp 1711653199
transform 1 0 2848 0 1 2570
box -8 -3 16 105
use FILL  FILL_571
timestamp 1711653199
transform 1 0 2840 0 1 2570
box -8 -3 16 105
use FILL  FILL_572
timestamp 1711653199
transform 1 0 2736 0 1 2570
box -8 -3 16 105
use FILL  FILL_573
timestamp 1711653199
transform 1 0 2728 0 1 2570
box -8 -3 16 105
use FILL  FILL_574
timestamp 1711653199
transform 1 0 2640 0 1 2570
box -8 -3 16 105
use FILL  FILL_575
timestamp 1711653199
transform 1 0 2536 0 1 2570
box -8 -3 16 105
use FILL  FILL_576
timestamp 1711653199
transform 1 0 2528 0 1 2570
box -8 -3 16 105
use FILL  FILL_577
timestamp 1711653199
transform 1 0 2424 0 1 2570
box -8 -3 16 105
use FILL  FILL_578
timestamp 1711653199
transform 1 0 2320 0 1 2570
box -8 -3 16 105
use FILL  FILL_579
timestamp 1711653199
transform 1 0 2216 0 1 2570
box -8 -3 16 105
use FILL  FILL_580
timestamp 1711653199
transform 1 0 2208 0 1 2570
box -8 -3 16 105
use FILL  FILL_581
timestamp 1711653199
transform 1 0 2200 0 1 2570
box -8 -3 16 105
use FILL  FILL_582
timestamp 1711653199
transform 1 0 2192 0 1 2570
box -8 -3 16 105
use FILL  FILL_583
timestamp 1711653199
transform 1 0 2104 0 1 2570
box -8 -3 16 105
use FILL  FILL_584
timestamp 1711653199
transform 1 0 2096 0 1 2570
box -8 -3 16 105
use FILL  FILL_585
timestamp 1711653199
transform 1 0 2088 0 1 2570
box -8 -3 16 105
use FILL  FILL_586
timestamp 1711653199
transform 1 0 2080 0 1 2570
box -8 -3 16 105
use FILL  FILL_587
timestamp 1711653199
transform 1 0 1984 0 1 2570
box -8 -3 16 105
use FILL  FILL_588
timestamp 1711653199
transform 1 0 1976 0 1 2570
box -8 -3 16 105
use FILL  FILL_589
timestamp 1711653199
transform 1 0 1968 0 1 2570
box -8 -3 16 105
use FILL  FILL_590
timestamp 1711653199
transform 1 0 1864 0 1 2570
box -8 -3 16 105
use FILL  FILL_591
timestamp 1711653199
transform 1 0 1824 0 1 2570
box -8 -3 16 105
use FILL  FILL_592
timestamp 1711653199
transform 1 0 1800 0 1 2570
box -8 -3 16 105
use FILL  FILL_593
timestamp 1711653199
transform 1 0 1696 0 1 2570
box -8 -3 16 105
use FILL  FILL_594
timestamp 1711653199
transform 1 0 1688 0 1 2570
box -8 -3 16 105
use FILL  FILL_595
timestamp 1711653199
transform 1 0 1680 0 1 2570
box -8 -3 16 105
use FILL  FILL_596
timestamp 1711653199
transform 1 0 1600 0 1 2570
box -8 -3 16 105
use FILL  FILL_597
timestamp 1711653199
transform 1 0 1592 0 1 2570
box -8 -3 16 105
use FILL  FILL_598
timestamp 1711653199
transform 1 0 1584 0 1 2570
box -8 -3 16 105
use FILL  FILL_599
timestamp 1711653199
transform 1 0 1480 0 1 2570
box -8 -3 16 105
use FILL  FILL_600
timestamp 1711653199
transform 1 0 1448 0 1 2570
box -8 -3 16 105
use FILL  FILL_601
timestamp 1711653199
transform 1 0 1344 0 1 2570
box -8 -3 16 105
use FILL  FILL_602
timestamp 1711653199
transform 1 0 1336 0 1 2570
box -8 -3 16 105
use FILL  FILL_603
timestamp 1711653199
transform 1 0 1328 0 1 2570
box -8 -3 16 105
use FILL  FILL_604
timestamp 1711653199
transform 1 0 1320 0 1 2570
box -8 -3 16 105
use FILL  FILL_605
timestamp 1711653199
transform 1 0 1256 0 1 2570
box -8 -3 16 105
use FILL  FILL_606
timestamp 1711653199
transform 1 0 1248 0 1 2570
box -8 -3 16 105
use FILL  FILL_607
timestamp 1711653199
transform 1 0 1240 0 1 2570
box -8 -3 16 105
use FILL  FILL_608
timestamp 1711653199
transform 1 0 1176 0 1 2570
box -8 -3 16 105
use FILL  FILL_609
timestamp 1711653199
transform 1 0 1168 0 1 2570
box -8 -3 16 105
use FILL  FILL_610
timestamp 1711653199
transform 1 0 1160 0 1 2570
box -8 -3 16 105
use FILL  FILL_611
timestamp 1711653199
transform 1 0 1088 0 1 2570
box -8 -3 16 105
use FILL  FILL_612
timestamp 1711653199
transform 1 0 1080 0 1 2570
box -8 -3 16 105
use FILL  FILL_613
timestamp 1711653199
transform 1 0 1048 0 1 2570
box -8 -3 16 105
use FILL  FILL_614
timestamp 1711653199
transform 1 0 1040 0 1 2570
box -8 -3 16 105
use FILL  FILL_615
timestamp 1711653199
transform 1 0 976 0 1 2570
box -8 -3 16 105
use FILL  FILL_616
timestamp 1711653199
transform 1 0 968 0 1 2570
box -8 -3 16 105
use FILL  FILL_617
timestamp 1711653199
transform 1 0 960 0 1 2570
box -8 -3 16 105
use FILL  FILL_618
timestamp 1711653199
transform 1 0 880 0 1 2570
box -8 -3 16 105
use FILL  FILL_619
timestamp 1711653199
transform 1 0 872 0 1 2570
box -8 -3 16 105
use FILL  FILL_620
timestamp 1711653199
transform 1 0 864 0 1 2570
box -8 -3 16 105
use FILL  FILL_621
timestamp 1711653199
transform 1 0 776 0 1 2570
box -8 -3 16 105
use FILL  FILL_622
timestamp 1711653199
transform 1 0 768 0 1 2570
box -8 -3 16 105
use FILL  FILL_623
timestamp 1711653199
transform 1 0 712 0 1 2570
box -8 -3 16 105
use FILL  FILL_624
timestamp 1711653199
transform 1 0 704 0 1 2570
box -8 -3 16 105
use FILL  FILL_625
timestamp 1711653199
transform 1 0 632 0 1 2570
box -8 -3 16 105
use FILL  FILL_626
timestamp 1711653199
transform 1 0 624 0 1 2570
box -8 -3 16 105
use FILL  FILL_627
timestamp 1711653199
transform 1 0 592 0 1 2570
box -8 -3 16 105
use FILL  FILL_628
timestamp 1711653199
transform 1 0 560 0 1 2570
box -8 -3 16 105
use FILL  FILL_629
timestamp 1711653199
transform 1 0 504 0 1 2570
box -8 -3 16 105
use FILL  FILL_630
timestamp 1711653199
transform 1 0 400 0 1 2570
box -8 -3 16 105
use FILL  FILL_631
timestamp 1711653199
transform 1 0 392 0 1 2570
box -8 -3 16 105
use FILL  FILL_632
timestamp 1711653199
transform 1 0 256 0 1 2570
box -8 -3 16 105
use FILL  FILL_633
timestamp 1711653199
transform 1 0 248 0 1 2570
box -8 -3 16 105
use FILL  FILL_634
timestamp 1711653199
transform 1 0 192 0 1 2570
box -8 -3 16 105
use FILL  FILL_635
timestamp 1711653199
transform 1 0 184 0 1 2570
box -8 -3 16 105
use FILL  FILL_636
timestamp 1711653199
transform 1 0 176 0 1 2570
box -8 -3 16 105
use FILL  FILL_637
timestamp 1711653199
transform 1 0 72 0 1 2570
box -8 -3 16 105
use FILL  FILL_638
timestamp 1711653199
transform 1 0 3392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_639
timestamp 1711653199
transform 1 0 3384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_640
timestamp 1711653199
transform 1 0 3312 0 -1 2570
box -8 -3 16 105
use FILL  FILL_641
timestamp 1711653199
transform 1 0 3304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_642
timestamp 1711653199
transform 1 0 3256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_643
timestamp 1711653199
transform 1 0 3248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_644
timestamp 1711653199
transform 1 0 3240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_645
timestamp 1711653199
transform 1 0 3184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_646
timestamp 1711653199
transform 1 0 3176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_647
timestamp 1711653199
transform 1 0 3168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_648
timestamp 1711653199
transform 1 0 3096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_649
timestamp 1711653199
transform 1 0 3088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_650
timestamp 1711653199
transform 1 0 2984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_651
timestamp 1711653199
transform 1 0 2976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_652
timestamp 1711653199
transform 1 0 2968 0 -1 2570
box -8 -3 16 105
use FILL  FILL_653
timestamp 1711653199
transform 1 0 2896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_654
timestamp 1711653199
transform 1 0 2792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_655
timestamp 1711653199
transform 1 0 2784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_656
timestamp 1711653199
transform 1 0 2776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_657
timestamp 1711653199
transform 1 0 2640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_658
timestamp 1711653199
transform 1 0 2536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_659
timestamp 1711653199
transform 1 0 2432 0 -1 2570
box -8 -3 16 105
use FILL  FILL_660
timestamp 1711653199
transform 1 0 2392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_661
timestamp 1711653199
transform 1 0 2384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_662
timestamp 1711653199
transform 1 0 2280 0 -1 2570
box -8 -3 16 105
use FILL  FILL_663
timestamp 1711653199
transform 1 0 2272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_664
timestamp 1711653199
transform 1 0 2168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_665
timestamp 1711653199
transform 1 0 2160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_666
timestamp 1711653199
transform 1 0 2152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_667
timestamp 1711653199
transform 1 0 2064 0 -1 2570
box -8 -3 16 105
use FILL  FILL_668
timestamp 1711653199
transform 1 0 2056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_669
timestamp 1711653199
transform 1 0 2048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_670
timestamp 1711653199
transform 1 0 1944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_671
timestamp 1711653199
transform 1 0 1840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_672
timestamp 1711653199
transform 1 0 1832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_673
timestamp 1711653199
transform 1 0 1824 0 -1 2570
box -8 -3 16 105
use FILL  FILL_674
timestamp 1711653199
transform 1 0 1736 0 -1 2570
box -8 -3 16 105
use FILL  FILL_675
timestamp 1711653199
transform 1 0 1728 0 -1 2570
box -8 -3 16 105
use FILL  FILL_676
timestamp 1711653199
transform 1 0 1720 0 -1 2570
box -8 -3 16 105
use FILL  FILL_677
timestamp 1711653199
transform 1 0 1712 0 -1 2570
box -8 -3 16 105
use FILL  FILL_678
timestamp 1711653199
transform 1 0 1624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_679
timestamp 1711653199
transform 1 0 1616 0 -1 2570
box -8 -3 16 105
use FILL  FILL_680
timestamp 1711653199
transform 1 0 1608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_681
timestamp 1711653199
transform 1 0 1600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_682
timestamp 1711653199
transform 1 0 1592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_683
timestamp 1711653199
transform 1 0 1520 0 -1 2570
box -8 -3 16 105
use FILL  FILL_684
timestamp 1711653199
transform 1 0 1512 0 -1 2570
box -8 -3 16 105
use FILL  FILL_685
timestamp 1711653199
transform 1 0 1456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_686
timestamp 1711653199
transform 1 0 1416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_687
timestamp 1711653199
transform 1 0 1360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_688
timestamp 1711653199
transform 1 0 1352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_689
timestamp 1711653199
transform 1 0 1248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_690
timestamp 1711653199
transform 1 0 1240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_691
timestamp 1711653199
transform 1 0 1232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_692
timestamp 1711653199
transform 1 0 1144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_693
timestamp 1711653199
transform 1 0 1136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_694
timestamp 1711653199
transform 1 0 1128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_695
timestamp 1711653199
transform 1 0 1080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_696
timestamp 1711653199
transform 1 0 1032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_697
timestamp 1711653199
transform 1 0 1024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_698
timestamp 1711653199
transform 1 0 984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_699
timestamp 1711653199
transform 1 0 976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_700
timestamp 1711653199
transform 1 0 968 0 -1 2570
box -8 -3 16 105
use FILL  FILL_701
timestamp 1711653199
transform 1 0 960 0 -1 2570
box -8 -3 16 105
use FILL  FILL_702
timestamp 1711653199
transform 1 0 880 0 -1 2570
box -8 -3 16 105
use FILL  FILL_703
timestamp 1711653199
transform 1 0 872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_704
timestamp 1711653199
transform 1 0 768 0 -1 2570
box -8 -3 16 105
use FILL  FILL_705
timestamp 1711653199
transform 1 0 760 0 -1 2570
box -8 -3 16 105
use FILL  FILL_706
timestamp 1711653199
transform 1 0 752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_707
timestamp 1711653199
transform 1 0 744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_708
timestamp 1711653199
transform 1 0 664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_709
timestamp 1711653199
transform 1 0 656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_710
timestamp 1711653199
transform 1 0 648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_711
timestamp 1711653199
transform 1 0 544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_712
timestamp 1711653199
transform 1 0 536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_713
timestamp 1711653199
transform 1 0 504 0 -1 2570
box -8 -3 16 105
use FILL  FILL_714
timestamp 1711653199
transform 1 0 400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_715
timestamp 1711653199
transform 1 0 392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_716
timestamp 1711653199
transform 1 0 384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_717
timestamp 1711653199
transform 1 0 376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_718
timestamp 1711653199
transform 1 0 368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_719
timestamp 1711653199
transform 1 0 320 0 -1 2570
box -8 -3 16 105
use FILL  FILL_720
timestamp 1711653199
transform 1 0 312 0 -1 2570
box -8 -3 16 105
use FILL  FILL_721
timestamp 1711653199
transform 1 0 304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_722
timestamp 1711653199
transform 1 0 296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_723
timestamp 1711653199
transform 1 0 288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_724
timestamp 1711653199
transform 1 0 280 0 -1 2570
box -8 -3 16 105
use FILL  FILL_725
timestamp 1711653199
transform 1 0 192 0 -1 2570
box -8 -3 16 105
use FILL  FILL_726
timestamp 1711653199
transform 1 0 184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_727
timestamp 1711653199
transform 1 0 176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_728
timestamp 1711653199
transform 1 0 72 0 -1 2570
box -8 -3 16 105
use FILL  FILL_729
timestamp 1711653199
transform 1 0 3392 0 1 2370
box -8 -3 16 105
use FILL  FILL_730
timestamp 1711653199
transform 1 0 3384 0 1 2370
box -8 -3 16 105
use FILL  FILL_731
timestamp 1711653199
transform 1 0 3376 0 1 2370
box -8 -3 16 105
use FILL  FILL_732
timestamp 1711653199
transform 1 0 3304 0 1 2370
box -8 -3 16 105
use FILL  FILL_733
timestamp 1711653199
transform 1 0 3296 0 1 2370
box -8 -3 16 105
use FILL  FILL_734
timestamp 1711653199
transform 1 0 3256 0 1 2370
box -8 -3 16 105
use FILL  FILL_735
timestamp 1711653199
transform 1 0 3248 0 1 2370
box -8 -3 16 105
use FILL  FILL_736
timestamp 1711653199
transform 1 0 3184 0 1 2370
box -8 -3 16 105
use FILL  FILL_737
timestamp 1711653199
transform 1 0 3176 0 1 2370
box -8 -3 16 105
use FILL  FILL_738
timestamp 1711653199
transform 1 0 3136 0 1 2370
box -8 -3 16 105
use FILL  FILL_739
timestamp 1711653199
transform 1 0 3096 0 1 2370
box -8 -3 16 105
use FILL  FILL_740
timestamp 1711653199
transform 1 0 3056 0 1 2370
box -8 -3 16 105
use FILL  FILL_741
timestamp 1711653199
transform 1 0 3048 0 1 2370
box -8 -3 16 105
use FILL  FILL_742
timestamp 1711653199
transform 1 0 3040 0 1 2370
box -8 -3 16 105
use FILL  FILL_743
timestamp 1711653199
transform 1 0 3032 0 1 2370
box -8 -3 16 105
use FILL  FILL_744
timestamp 1711653199
transform 1 0 2824 0 1 2370
box -8 -3 16 105
use FILL  FILL_745
timestamp 1711653199
transform 1 0 2816 0 1 2370
box -8 -3 16 105
use FILL  FILL_746
timestamp 1711653199
transform 1 0 2728 0 1 2370
box -8 -3 16 105
use FILL  FILL_747
timestamp 1711653199
transform 1 0 2624 0 1 2370
box -8 -3 16 105
use FILL  FILL_748
timestamp 1711653199
transform 1 0 2616 0 1 2370
box -8 -3 16 105
use FILL  FILL_749
timestamp 1711653199
transform 1 0 2480 0 1 2370
box -8 -3 16 105
use FILL  FILL_750
timestamp 1711653199
transform 1 0 2472 0 1 2370
box -8 -3 16 105
use FILL  FILL_751
timestamp 1711653199
transform 1 0 2400 0 1 2370
box -8 -3 16 105
use FILL  FILL_752
timestamp 1711653199
transform 1 0 2392 0 1 2370
box -8 -3 16 105
use FILL  FILL_753
timestamp 1711653199
transform 1 0 2352 0 1 2370
box -8 -3 16 105
use FILL  FILL_754
timestamp 1711653199
transform 1 0 2312 0 1 2370
box -8 -3 16 105
use FILL  FILL_755
timestamp 1711653199
transform 1 0 2304 0 1 2370
box -8 -3 16 105
use FILL  FILL_756
timestamp 1711653199
transform 1 0 2232 0 1 2370
box -8 -3 16 105
use FILL  FILL_757
timestamp 1711653199
transform 1 0 2224 0 1 2370
box -8 -3 16 105
use FILL  FILL_758
timestamp 1711653199
transform 1 0 2120 0 1 2370
box -8 -3 16 105
use FILL  FILL_759
timestamp 1711653199
transform 1 0 2016 0 1 2370
box -8 -3 16 105
use FILL  FILL_760
timestamp 1711653199
transform 1 0 1872 0 1 2370
box -8 -3 16 105
use FILL  FILL_761
timestamp 1711653199
transform 1 0 1864 0 1 2370
box -8 -3 16 105
use FILL  FILL_762
timestamp 1711653199
transform 1 0 1760 0 1 2370
box -8 -3 16 105
use FILL  FILL_763
timestamp 1711653199
transform 1 0 1752 0 1 2370
box -8 -3 16 105
use FILL  FILL_764
timestamp 1711653199
transform 1 0 1744 0 1 2370
box -8 -3 16 105
use FILL  FILL_765
timestamp 1711653199
transform 1 0 1664 0 1 2370
box -8 -3 16 105
use FILL  FILL_766
timestamp 1711653199
transform 1 0 1640 0 1 2370
box -8 -3 16 105
use FILL  FILL_767
timestamp 1711653199
transform 1 0 1592 0 1 2370
box -8 -3 16 105
use FILL  FILL_768
timestamp 1711653199
transform 1 0 1488 0 1 2370
box -8 -3 16 105
use FILL  FILL_769
timestamp 1711653199
transform 1 0 1480 0 1 2370
box -8 -3 16 105
use FILL  FILL_770
timestamp 1711653199
transform 1 0 1472 0 1 2370
box -8 -3 16 105
use FILL  FILL_771
timestamp 1711653199
transform 1 0 1376 0 1 2370
box -8 -3 16 105
use FILL  FILL_772
timestamp 1711653199
transform 1 0 1368 0 1 2370
box -8 -3 16 105
use FILL  FILL_773
timestamp 1711653199
transform 1 0 1360 0 1 2370
box -8 -3 16 105
use FILL  FILL_774
timestamp 1711653199
transform 1 0 1352 0 1 2370
box -8 -3 16 105
use FILL  FILL_775
timestamp 1711653199
transform 1 0 1344 0 1 2370
box -8 -3 16 105
use FILL  FILL_776
timestamp 1711653199
transform 1 0 1264 0 1 2370
box -8 -3 16 105
use FILL  FILL_777
timestamp 1711653199
transform 1 0 1256 0 1 2370
box -8 -3 16 105
use FILL  FILL_778
timestamp 1711653199
transform 1 0 1248 0 1 2370
box -8 -3 16 105
use FILL  FILL_779
timestamp 1711653199
transform 1 0 1176 0 1 2370
box -8 -3 16 105
use FILL  FILL_780
timestamp 1711653199
transform 1 0 1168 0 1 2370
box -8 -3 16 105
use FILL  FILL_781
timestamp 1711653199
transform 1 0 1160 0 1 2370
box -8 -3 16 105
use FILL  FILL_782
timestamp 1711653199
transform 1 0 1072 0 1 2370
box -8 -3 16 105
use FILL  FILL_783
timestamp 1711653199
transform 1 0 1064 0 1 2370
box -8 -3 16 105
use FILL  FILL_784
timestamp 1711653199
transform 1 0 960 0 1 2370
box -8 -3 16 105
use FILL  FILL_785
timestamp 1711653199
transform 1 0 928 0 1 2370
box -8 -3 16 105
use FILL  FILL_786
timestamp 1711653199
transform 1 0 824 0 1 2370
box -8 -3 16 105
use FILL  FILL_787
timestamp 1711653199
transform 1 0 816 0 1 2370
box -8 -3 16 105
use FILL  FILL_788
timestamp 1711653199
transform 1 0 712 0 1 2370
box -8 -3 16 105
use FILL  FILL_789
timestamp 1711653199
transform 1 0 680 0 1 2370
box -8 -3 16 105
use FILL  FILL_790
timestamp 1711653199
transform 1 0 672 0 1 2370
box -8 -3 16 105
use FILL  FILL_791
timestamp 1711653199
transform 1 0 664 0 1 2370
box -8 -3 16 105
use FILL  FILL_792
timestamp 1711653199
transform 1 0 560 0 1 2370
box -8 -3 16 105
use FILL  FILL_793
timestamp 1711653199
transform 1 0 552 0 1 2370
box -8 -3 16 105
use FILL  FILL_794
timestamp 1711653199
transform 1 0 544 0 1 2370
box -8 -3 16 105
use FILL  FILL_795
timestamp 1711653199
transform 1 0 440 0 1 2370
box -8 -3 16 105
use FILL  FILL_796
timestamp 1711653199
transform 1 0 432 0 1 2370
box -8 -3 16 105
use FILL  FILL_797
timestamp 1711653199
transform 1 0 424 0 1 2370
box -8 -3 16 105
use FILL  FILL_798
timestamp 1711653199
transform 1 0 320 0 1 2370
box -8 -3 16 105
use FILL  FILL_799
timestamp 1711653199
transform 1 0 312 0 1 2370
box -8 -3 16 105
use FILL  FILL_800
timestamp 1711653199
transform 1 0 304 0 1 2370
box -8 -3 16 105
use FILL  FILL_801
timestamp 1711653199
transform 1 0 296 0 1 2370
box -8 -3 16 105
use FILL  FILL_802
timestamp 1711653199
transform 1 0 288 0 1 2370
box -8 -3 16 105
use FILL  FILL_803
timestamp 1711653199
transform 1 0 280 0 1 2370
box -8 -3 16 105
use FILL  FILL_804
timestamp 1711653199
transform 1 0 272 0 1 2370
box -8 -3 16 105
use FILL  FILL_805
timestamp 1711653199
transform 1 0 264 0 1 2370
box -8 -3 16 105
use FILL  FILL_806
timestamp 1711653199
transform 1 0 256 0 1 2370
box -8 -3 16 105
use FILL  FILL_807
timestamp 1711653199
transform 1 0 248 0 1 2370
box -8 -3 16 105
use FILL  FILL_808
timestamp 1711653199
transform 1 0 240 0 1 2370
box -8 -3 16 105
use FILL  FILL_809
timestamp 1711653199
transform 1 0 232 0 1 2370
box -8 -3 16 105
use FILL  FILL_810
timestamp 1711653199
transform 1 0 224 0 1 2370
box -8 -3 16 105
use FILL  FILL_811
timestamp 1711653199
transform 1 0 216 0 1 2370
box -8 -3 16 105
use FILL  FILL_812
timestamp 1711653199
transform 1 0 208 0 1 2370
box -8 -3 16 105
use FILL  FILL_813
timestamp 1711653199
transform 1 0 200 0 1 2370
box -8 -3 16 105
use FILL  FILL_814
timestamp 1711653199
transform 1 0 192 0 1 2370
box -8 -3 16 105
use FILL  FILL_815
timestamp 1711653199
transform 1 0 184 0 1 2370
box -8 -3 16 105
use FILL  FILL_816
timestamp 1711653199
transform 1 0 176 0 1 2370
box -8 -3 16 105
use FILL  FILL_817
timestamp 1711653199
transform 1 0 168 0 1 2370
box -8 -3 16 105
use FILL  FILL_818
timestamp 1711653199
transform 1 0 160 0 1 2370
box -8 -3 16 105
use FILL  FILL_819
timestamp 1711653199
transform 1 0 152 0 1 2370
box -8 -3 16 105
use FILL  FILL_820
timestamp 1711653199
transform 1 0 144 0 1 2370
box -8 -3 16 105
use FILL  FILL_821
timestamp 1711653199
transform 1 0 136 0 1 2370
box -8 -3 16 105
use FILL  FILL_822
timestamp 1711653199
transform 1 0 128 0 1 2370
box -8 -3 16 105
use FILL  FILL_823
timestamp 1711653199
transform 1 0 120 0 1 2370
box -8 -3 16 105
use FILL  FILL_824
timestamp 1711653199
transform 1 0 112 0 1 2370
box -8 -3 16 105
use FILL  FILL_825
timestamp 1711653199
transform 1 0 104 0 1 2370
box -8 -3 16 105
use FILL  FILL_826
timestamp 1711653199
transform 1 0 96 0 1 2370
box -8 -3 16 105
use FILL  FILL_827
timestamp 1711653199
transform 1 0 88 0 1 2370
box -8 -3 16 105
use FILL  FILL_828
timestamp 1711653199
transform 1 0 80 0 1 2370
box -8 -3 16 105
use FILL  FILL_829
timestamp 1711653199
transform 1 0 72 0 1 2370
box -8 -3 16 105
use FILL  FILL_830
timestamp 1711653199
transform 1 0 3392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_831
timestamp 1711653199
transform 1 0 3384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_832
timestamp 1711653199
transform 1 0 3376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_833
timestamp 1711653199
transform 1 0 3304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_834
timestamp 1711653199
transform 1 0 3296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_835
timestamp 1711653199
transform 1 0 3288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_836
timestamp 1711653199
transform 1 0 3280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_837
timestamp 1711653199
transform 1 0 3272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_838
timestamp 1711653199
transform 1 0 3200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_839
timestamp 1711653199
transform 1 0 3192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_840
timestamp 1711653199
transform 1 0 3184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_841
timestamp 1711653199
transform 1 0 3176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_842
timestamp 1711653199
transform 1 0 3168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_843
timestamp 1711653199
transform 1 0 3104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_844
timestamp 1711653199
transform 1 0 3096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_845
timestamp 1711653199
transform 1 0 3088 0 -1 2370
box -8 -3 16 105
use FILL  FILL_846
timestamp 1711653199
transform 1 0 2984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_847
timestamp 1711653199
transform 1 0 2976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_848
timestamp 1711653199
transform 1 0 2904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_849
timestamp 1711653199
transform 1 0 2896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_850
timestamp 1711653199
transform 1 0 2888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_851
timestamp 1711653199
transform 1 0 2880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_852
timestamp 1711653199
transform 1 0 2872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_853
timestamp 1711653199
transform 1 0 2832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_854
timestamp 1711653199
transform 1 0 2784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_855
timestamp 1711653199
transform 1 0 2776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_856
timestamp 1711653199
transform 1 0 2768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_857
timestamp 1711653199
transform 1 0 2760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_858
timestamp 1711653199
transform 1 0 2752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_859
timestamp 1711653199
transform 1 0 2696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_860
timestamp 1711653199
transform 1 0 2688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_861
timestamp 1711653199
transform 1 0 2680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_862
timestamp 1711653199
transform 1 0 2576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_863
timestamp 1711653199
transform 1 0 2568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_864
timestamp 1711653199
transform 1 0 2560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_865
timestamp 1711653199
transform 1 0 2552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_866
timestamp 1711653199
transform 1 0 2448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_867
timestamp 1711653199
transform 1 0 2440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_868
timestamp 1711653199
transform 1 0 2432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_869
timestamp 1711653199
transform 1 0 2360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_870
timestamp 1711653199
transform 1 0 2352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_871
timestamp 1711653199
transform 1 0 2344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_872
timestamp 1711653199
transform 1 0 2336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_873
timestamp 1711653199
transform 1 0 2328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_874
timestamp 1711653199
transform 1 0 2320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_875
timestamp 1711653199
transform 1 0 2264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_876
timestamp 1711653199
transform 1 0 2256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_877
timestamp 1711653199
transform 1 0 2232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_878
timestamp 1711653199
transform 1 0 2224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_879
timestamp 1711653199
transform 1 0 2216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_880
timestamp 1711653199
transform 1 0 2208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_881
timestamp 1711653199
transform 1 0 2144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_882
timestamp 1711653199
transform 1 0 2136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_883
timestamp 1711653199
transform 1 0 2128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_884
timestamp 1711653199
transform 1 0 2120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_885
timestamp 1711653199
transform 1 0 2096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_886
timestamp 1711653199
transform 1 0 2056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_887
timestamp 1711653199
transform 1 0 2048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_888
timestamp 1711653199
transform 1 0 2040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_889
timestamp 1711653199
transform 1 0 2032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_890
timestamp 1711653199
transform 1 0 1992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_891
timestamp 1711653199
transform 1 0 1984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_892
timestamp 1711653199
transform 1 0 1960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_893
timestamp 1711653199
transform 1 0 1952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_894
timestamp 1711653199
transform 1 0 1944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_895
timestamp 1711653199
transform 1 0 1936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_896
timestamp 1711653199
transform 1 0 1896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_897
timestamp 1711653199
transform 1 0 1888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_898
timestamp 1711653199
transform 1 0 1880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_899
timestamp 1711653199
transform 1 0 1872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_900
timestamp 1711653199
transform 1 0 1768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_901
timestamp 1711653199
transform 1 0 1760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_902
timestamp 1711653199
transform 1 0 1752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_903
timestamp 1711653199
transform 1 0 1744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_904
timestamp 1711653199
transform 1 0 1704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_905
timestamp 1711653199
transform 1 0 1696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_906
timestamp 1711653199
transform 1 0 1688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_907
timestamp 1711653199
transform 1 0 1616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_908
timestamp 1711653199
transform 1 0 1608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_909
timestamp 1711653199
transform 1 0 1600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_910
timestamp 1711653199
transform 1 0 1496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_911
timestamp 1711653199
transform 1 0 1488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_912
timestamp 1711653199
transform 1 0 1480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_913
timestamp 1711653199
transform 1 0 1440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_914
timestamp 1711653199
transform 1 0 1336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_915
timestamp 1711653199
transform 1 0 1328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_916
timestamp 1711653199
transform 1 0 1320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_917
timestamp 1711653199
transform 1 0 1312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_918
timestamp 1711653199
transform 1 0 1304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_919
timestamp 1711653199
transform 1 0 1264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_920
timestamp 1711653199
transform 1 0 1256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_921
timestamp 1711653199
transform 1 0 1248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_922
timestamp 1711653199
transform 1 0 1240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_923
timestamp 1711653199
transform 1 0 1136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_924
timestamp 1711653199
transform 1 0 1128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_925
timestamp 1711653199
transform 1 0 1024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_926
timestamp 1711653199
transform 1 0 1016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_927
timestamp 1711653199
transform 1 0 1008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_928
timestamp 1711653199
transform 1 0 1000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_929
timestamp 1711653199
transform 1 0 992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_930
timestamp 1711653199
transform 1 0 984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_931
timestamp 1711653199
transform 1 0 912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_932
timestamp 1711653199
transform 1 0 904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_933
timestamp 1711653199
transform 1 0 896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_934
timestamp 1711653199
transform 1 0 792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_935
timestamp 1711653199
transform 1 0 784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_936
timestamp 1711653199
transform 1 0 776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_937
timestamp 1711653199
transform 1 0 672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_938
timestamp 1711653199
transform 1 0 664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_939
timestamp 1711653199
transform 1 0 656 0 -1 2370
box -8 -3 16 105
use FILL  FILL_940
timestamp 1711653199
transform 1 0 616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_941
timestamp 1711653199
transform 1 0 608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_942
timestamp 1711653199
transform 1 0 504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_943
timestamp 1711653199
transform 1 0 496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_944
timestamp 1711653199
transform 1 0 392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_945
timestamp 1711653199
transform 1 0 288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_946
timestamp 1711653199
transform 1 0 280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_947
timestamp 1711653199
transform 1 0 176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_948
timestamp 1711653199
transform 1 0 72 0 -1 2370
box -8 -3 16 105
use FILL  FILL_949
timestamp 1711653199
transform 1 0 3392 0 1 2170
box -8 -3 16 105
use FILL  FILL_950
timestamp 1711653199
transform 1 0 3384 0 1 2170
box -8 -3 16 105
use FILL  FILL_951
timestamp 1711653199
transform 1 0 3288 0 1 2170
box -8 -3 16 105
use FILL  FILL_952
timestamp 1711653199
transform 1 0 3280 0 1 2170
box -8 -3 16 105
use FILL  FILL_953
timestamp 1711653199
transform 1 0 3272 0 1 2170
box -8 -3 16 105
use FILL  FILL_954
timestamp 1711653199
transform 1 0 3264 0 1 2170
box -8 -3 16 105
use FILL  FILL_955
timestamp 1711653199
transform 1 0 3256 0 1 2170
box -8 -3 16 105
use FILL  FILL_956
timestamp 1711653199
transform 1 0 3248 0 1 2170
box -8 -3 16 105
use FILL  FILL_957
timestamp 1711653199
transform 1 0 3184 0 1 2170
box -8 -3 16 105
use FILL  FILL_958
timestamp 1711653199
transform 1 0 3176 0 1 2170
box -8 -3 16 105
use FILL  FILL_959
timestamp 1711653199
transform 1 0 3168 0 1 2170
box -8 -3 16 105
use FILL  FILL_960
timestamp 1711653199
transform 1 0 3136 0 1 2170
box -8 -3 16 105
use FILL  FILL_961
timestamp 1711653199
transform 1 0 3080 0 1 2170
box -8 -3 16 105
use FILL  FILL_962
timestamp 1711653199
transform 1 0 3072 0 1 2170
box -8 -3 16 105
use FILL  FILL_963
timestamp 1711653199
transform 1 0 3064 0 1 2170
box -8 -3 16 105
use FILL  FILL_964
timestamp 1711653199
transform 1 0 2960 0 1 2170
box -8 -3 16 105
use FILL  FILL_965
timestamp 1711653199
transform 1 0 2856 0 1 2170
box -8 -3 16 105
use FILL  FILL_966
timestamp 1711653199
transform 1 0 2848 0 1 2170
box -8 -3 16 105
use FILL  FILL_967
timestamp 1711653199
transform 1 0 2744 0 1 2170
box -8 -3 16 105
use FILL  FILL_968
timestamp 1711653199
transform 1 0 2736 0 1 2170
box -8 -3 16 105
use FILL  FILL_969
timestamp 1711653199
transform 1 0 2544 0 1 2170
box -8 -3 16 105
use FILL  FILL_970
timestamp 1711653199
transform 1 0 2472 0 1 2170
box -8 -3 16 105
use FILL  FILL_971
timestamp 1711653199
transform 1 0 2464 0 1 2170
box -8 -3 16 105
use FILL  FILL_972
timestamp 1711653199
transform 1 0 2456 0 1 2170
box -8 -3 16 105
use FILL  FILL_973
timestamp 1711653199
transform 1 0 2416 0 1 2170
box -8 -3 16 105
use FILL  FILL_974
timestamp 1711653199
transform 1 0 2344 0 1 2170
box -8 -3 16 105
use FILL  FILL_975
timestamp 1711653199
transform 1 0 2336 0 1 2170
box -8 -3 16 105
use FILL  FILL_976
timestamp 1711653199
transform 1 0 2264 0 1 2170
box -8 -3 16 105
use FILL  FILL_977
timestamp 1711653199
transform 1 0 2256 0 1 2170
box -8 -3 16 105
use FILL  FILL_978
timestamp 1711653199
transform 1 0 2184 0 1 2170
box -8 -3 16 105
use FILL  FILL_979
timestamp 1711653199
transform 1 0 2160 0 1 2170
box -8 -3 16 105
use FILL  FILL_980
timestamp 1711653199
transform 1 0 2152 0 1 2170
box -8 -3 16 105
use FILL  FILL_981
timestamp 1711653199
transform 1 0 2144 0 1 2170
box -8 -3 16 105
use FILL  FILL_982
timestamp 1711653199
transform 1 0 2048 0 1 2170
box -8 -3 16 105
use FILL  FILL_983
timestamp 1711653199
transform 1 0 2040 0 1 2170
box -8 -3 16 105
use FILL  FILL_984
timestamp 1711653199
transform 1 0 2000 0 1 2170
box -8 -3 16 105
use FILL  FILL_985
timestamp 1711653199
transform 1 0 1992 0 1 2170
box -8 -3 16 105
use FILL  FILL_986
timestamp 1711653199
transform 1 0 1960 0 1 2170
box -8 -3 16 105
use FILL  FILL_987
timestamp 1711653199
transform 1 0 1920 0 1 2170
box -8 -3 16 105
use FILL  FILL_988
timestamp 1711653199
transform 1 0 1896 0 1 2170
box -8 -3 16 105
use FILL  FILL_989
timestamp 1711653199
transform 1 0 1848 0 1 2170
box -8 -3 16 105
use FILL  FILL_990
timestamp 1711653199
transform 1 0 1808 0 1 2170
box -8 -3 16 105
use FILL  FILL_991
timestamp 1711653199
transform 1 0 1768 0 1 2170
box -8 -3 16 105
use FILL  FILL_992
timestamp 1711653199
transform 1 0 1760 0 1 2170
box -8 -3 16 105
use FILL  FILL_993
timestamp 1711653199
transform 1 0 1720 0 1 2170
box -8 -3 16 105
use FILL  FILL_994
timestamp 1711653199
transform 1 0 1712 0 1 2170
box -8 -3 16 105
use FILL  FILL_995
timestamp 1711653199
transform 1 0 1704 0 1 2170
box -8 -3 16 105
use FILL  FILL_996
timestamp 1711653199
transform 1 0 1696 0 1 2170
box -8 -3 16 105
use FILL  FILL_997
timestamp 1711653199
transform 1 0 1688 0 1 2170
box -8 -3 16 105
use FILL  FILL_998
timestamp 1711653199
transform 1 0 1648 0 1 2170
box -8 -3 16 105
use FILL  FILL_999
timestamp 1711653199
transform 1 0 1640 0 1 2170
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1711653199
transform 1 0 1608 0 1 2170
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1711653199
transform 1 0 1600 0 1 2170
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1711653199
transform 1 0 1592 0 1 2170
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1711653199
transform 1 0 1584 0 1 2170
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1711653199
transform 1 0 1552 0 1 2170
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1711653199
transform 1 0 1544 0 1 2170
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1711653199
transform 1 0 1536 0 1 2170
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1711653199
transform 1 0 1488 0 1 2170
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1711653199
transform 1 0 1480 0 1 2170
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1711653199
transform 1 0 1472 0 1 2170
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1711653199
transform 1 0 1464 0 1 2170
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1711653199
transform 1 0 1432 0 1 2170
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1711653199
transform 1 0 1424 0 1 2170
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1711653199
transform 1 0 1416 0 1 2170
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1711653199
transform 1 0 1376 0 1 2170
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1711653199
transform 1 0 1368 0 1 2170
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1711653199
transform 1 0 1360 0 1 2170
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1711653199
transform 1 0 1352 0 1 2170
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1711653199
transform 1 0 1344 0 1 2170
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1711653199
transform 1 0 1320 0 1 2170
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1711653199
transform 1 0 1288 0 1 2170
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1711653199
transform 1 0 1280 0 1 2170
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1711653199
transform 1 0 1272 0 1 2170
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1711653199
transform 1 0 1264 0 1 2170
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1711653199
transform 1 0 1256 0 1 2170
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1711653199
transform 1 0 1216 0 1 2170
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1711653199
transform 1 0 1208 0 1 2170
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1711653199
transform 1 0 1200 0 1 2170
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1711653199
transform 1 0 1168 0 1 2170
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1711653199
transform 1 0 1160 0 1 2170
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1711653199
transform 1 0 1104 0 1 2170
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1711653199
transform 1 0 1096 0 1 2170
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1711653199
transform 1 0 1064 0 1 2170
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1711653199
transform 1 0 1056 0 1 2170
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1711653199
transform 1 0 1048 0 1 2170
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1711653199
transform 1 0 1040 0 1 2170
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1711653199
transform 1 0 1032 0 1 2170
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1711653199
transform 1 0 992 0 1 2170
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1711653199
transform 1 0 984 0 1 2170
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1711653199
transform 1 0 976 0 1 2170
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1711653199
transform 1 0 968 0 1 2170
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1711653199
transform 1 0 960 0 1 2170
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1711653199
transform 1 0 920 0 1 2170
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1711653199
transform 1 0 912 0 1 2170
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1711653199
transform 1 0 904 0 1 2170
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1711653199
transform 1 0 896 0 1 2170
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1711653199
transform 1 0 888 0 1 2170
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1711653199
transform 1 0 840 0 1 2170
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1711653199
transform 1 0 832 0 1 2170
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1711653199
transform 1 0 824 0 1 2170
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1711653199
transform 1 0 816 0 1 2170
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1711653199
transform 1 0 808 0 1 2170
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1711653199
transform 1 0 760 0 1 2170
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1711653199
transform 1 0 752 0 1 2170
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1711653199
transform 1 0 728 0 1 2170
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1711653199
transform 1 0 720 0 1 2170
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1711653199
transform 1 0 712 0 1 2170
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1711653199
transform 1 0 704 0 1 2170
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1711653199
transform 1 0 696 0 1 2170
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1711653199
transform 1 0 688 0 1 2170
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1711653199
transform 1 0 640 0 1 2170
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1711653199
transform 1 0 616 0 1 2170
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1711653199
transform 1 0 608 0 1 2170
box -8 -3 16 105
use FILL  FILL_1063
timestamp 1711653199
transform 1 0 600 0 1 2170
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1711653199
transform 1 0 592 0 1 2170
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1711653199
transform 1 0 520 0 1 2170
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1711653199
transform 1 0 512 0 1 2170
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1711653199
transform 1 0 472 0 1 2170
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1711653199
transform 1 0 464 0 1 2170
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1711653199
transform 1 0 456 0 1 2170
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1711653199
transform 1 0 448 0 1 2170
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1711653199
transform 1 0 392 0 1 2170
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1711653199
transform 1 0 384 0 1 2170
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1711653199
transform 1 0 376 0 1 2170
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1711653199
transform 1 0 368 0 1 2170
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1711653199
transform 1 0 312 0 1 2170
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1711653199
transform 1 0 304 0 1 2170
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1711653199
transform 1 0 296 0 1 2170
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1711653199
transform 1 0 288 0 1 2170
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1711653199
transform 1 0 280 0 1 2170
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1711653199
transform 1 0 192 0 1 2170
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1711653199
transform 1 0 184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1711653199
transform 1 0 176 0 1 2170
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1711653199
transform 1 0 72 0 1 2170
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1711653199
transform 1 0 3392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1711653199
transform 1 0 3384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1711653199
transform 1 0 3376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1711653199
transform 1 0 3280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1711653199
transform 1 0 3176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1711653199
transform 1 0 3168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1711653199
transform 1 0 3080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1711653199
transform 1 0 3072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1711653199
transform 1 0 3064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1711653199
transform 1 0 2960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1711653199
transform 1 0 2952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1711653199
transform 1 0 2944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1711653199
transform 1 0 2936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1711653199
transform 1 0 2872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1711653199
transform 1 0 2808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1711653199
transform 1 0 2800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1711653199
transform 1 0 2792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1711653199
transform 1 0 2784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1711653199
transform 1 0 2744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1711653199
transform 1 0 2720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1711653199
transform 1 0 2712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1711653199
transform 1 0 2704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1711653199
transform 1 0 2664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1711653199
transform 1 0 2656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1711653199
transform 1 0 2648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1711653199
transform 1 0 2640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1711653199
transform 1 0 2600 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1711653199
transform 1 0 2560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1711653199
transform 1 0 2552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1711653199
transform 1 0 2544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1711653199
transform 1 0 2488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1711653199
transform 1 0 2480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1711653199
transform 1 0 2472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1711653199
transform 1 0 2464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1711653199
transform 1 0 2400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1711653199
transform 1 0 2376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1711653199
transform 1 0 2344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1711653199
transform 1 0 2336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1711653199
transform 1 0 2288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1711653199
transform 1 0 2280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1711653199
transform 1 0 2272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1711653199
transform 1 0 2264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1711653199
transform 1 0 2256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1711653199
transform 1 0 2200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1711653199
transform 1 0 2144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1711653199
transform 1 0 2136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1711653199
transform 1 0 2128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1711653199
transform 1 0 2120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1711653199
transform 1 0 2080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1711653199
transform 1 0 2032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1711653199
transform 1 0 2024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1711653199
transform 1 0 2016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1711653199
transform 1 0 2008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1711653199
transform 1 0 2000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1711653199
transform 1 0 1920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1711653199
transform 1 0 1912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1711653199
transform 1 0 1904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1711653199
transform 1 0 1824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1711653199
transform 1 0 1816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1711653199
transform 1 0 1808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1711653199
transform 1 0 1760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1711653199
transform 1 0 1720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1146
timestamp 1711653199
transform 1 0 1680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1711653199
transform 1 0 1672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1711653199
transform 1 0 1632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1711653199
transform 1 0 1624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1711653199
transform 1 0 1616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1711653199
transform 1 0 1568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1711653199
transform 1 0 1560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1711653199
transform 1 0 1552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1711653199
transform 1 0 1544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1711653199
transform 1 0 1536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1711653199
transform 1 0 1528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1711653199
transform 1 0 1480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1711653199
transform 1 0 1472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1711653199
transform 1 0 1464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1711653199
transform 1 0 1456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1711653199
transform 1 0 1416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1711653199
transform 1 0 1408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1711653199
transform 1 0 1400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1711653199
transform 1 0 1392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1711653199
transform 1 0 1384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1711653199
transform 1 0 1344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1167
timestamp 1711653199
transform 1 0 1336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1711653199
transform 1 0 1328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1711653199
transform 1 0 1320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1711653199
transform 1 0 1312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1711653199
transform 1 0 1272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1711653199
transform 1 0 1264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1711653199
transform 1 0 1232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1711653199
transform 1 0 1224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1711653199
transform 1 0 1216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1711653199
transform 1 0 1208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1711653199
transform 1 0 1160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1711653199
transform 1 0 1152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1711653199
transform 1 0 1144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1711653199
transform 1 0 1136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1711653199
transform 1 0 1112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1711653199
transform 1 0 1104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1711653199
transform 1 0 1064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1184
timestamp 1711653199
transform 1 0 1056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1711653199
transform 1 0 1048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1711653199
transform 1 0 1040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1711653199
transform 1 0 1000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1711653199
transform 1 0 992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1711653199
transform 1 0 984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1711653199
transform 1 0 976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1711653199
transform 1 0 928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1711653199
transform 1 0 920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1711653199
transform 1 0 912 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1711653199
transform 1 0 840 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1711653199
transform 1 0 832 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1711653199
transform 1 0 824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1711653199
transform 1 0 816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1711653199
transform 1 0 808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1711653199
transform 1 0 744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1711653199
transform 1 0 736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1711653199
transform 1 0 728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1202
timestamp 1711653199
transform 1 0 720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1711653199
transform 1 0 712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1711653199
transform 1 0 688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1711653199
transform 1 0 640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1711653199
transform 1 0 632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1711653199
transform 1 0 624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1711653199
transform 1 0 560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1711653199
transform 1 0 552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1711653199
transform 1 0 512 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1711653199
transform 1 0 504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1711653199
transform 1 0 440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1711653199
transform 1 0 432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1711653199
transform 1 0 424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1711653199
transform 1 0 384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1711653199
transform 1 0 344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1217
timestamp 1711653199
transform 1 0 336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1711653199
transform 1 0 304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1711653199
transform 1 0 296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1711653199
transform 1 0 224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1221
timestamp 1711653199
transform 1 0 216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1711653199
transform 1 0 152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1711653199
transform 1 0 144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1711653199
transform 1 0 136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1711653199
transform 1 0 128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1711653199
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1711653199
transform 1 0 3392 0 1 1970
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1711653199
transform 1 0 3384 0 1 1970
box -8 -3 16 105
use FILL  FILL_1229
timestamp 1711653199
transform 1 0 3376 0 1 1970
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1711653199
transform 1 0 3368 0 1 1970
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1711653199
transform 1 0 3360 0 1 1970
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1711653199
transform 1 0 3352 0 1 1970
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1711653199
transform 1 0 3248 0 1 1970
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1711653199
transform 1 0 3240 0 1 1970
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1711653199
transform 1 0 3232 0 1 1970
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1711653199
transform 1 0 3224 0 1 1970
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1711653199
transform 1 0 3216 0 1 1970
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1711653199
transform 1 0 3208 0 1 1970
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1711653199
transform 1 0 3200 0 1 1970
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1711653199
transform 1 0 3192 0 1 1970
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1711653199
transform 1 0 3184 0 1 1970
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1711653199
transform 1 0 3176 0 1 1970
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1711653199
transform 1 0 3168 0 1 1970
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1711653199
transform 1 0 3160 0 1 1970
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1711653199
transform 1 0 3120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1711653199
transform 1 0 3112 0 1 1970
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1711653199
transform 1 0 3104 0 1 1970
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1711653199
transform 1 0 3096 0 1 1970
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1711653199
transform 1 0 3088 0 1 1970
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1711653199
transform 1 0 3048 0 1 1970
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1711653199
transform 1 0 3040 0 1 1970
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1711653199
transform 1 0 3032 0 1 1970
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1711653199
transform 1 0 2992 0 1 1970
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1711653199
transform 1 0 2984 0 1 1970
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1711653199
transform 1 0 2976 0 1 1970
box -8 -3 16 105
use FILL  FILL_1256
timestamp 1711653199
transform 1 0 2968 0 1 1970
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1711653199
transform 1 0 2944 0 1 1970
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1711653199
transform 1 0 2936 0 1 1970
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1711653199
transform 1 0 2896 0 1 1970
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1711653199
transform 1 0 2888 0 1 1970
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1711653199
transform 1 0 2880 0 1 1970
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1711653199
transform 1 0 2832 0 1 1970
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1711653199
transform 1 0 2824 0 1 1970
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1711653199
transform 1 0 2816 0 1 1970
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1711653199
transform 1 0 2776 0 1 1970
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1711653199
transform 1 0 2768 0 1 1970
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1711653199
transform 1 0 2720 0 1 1970
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1711653199
transform 1 0 2712 0 1 1970
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1711653199
transform 1 0 2704 0 1 1970
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1711653199
transform 1 0 2696 0 1 1970
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1711653199
transform 1 0 2656 0 1 1970
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1711653199
transform 1 0 2608 0 1 1970
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1711653199
transform 1 0 2600 0 1 1970
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1711653199
transform 1 0 2592 0 1 1970
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1711653199
transform 1 0 2584 0 1 1970
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1711653199
transform 1 0 2576 0 1 1970
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1711653199
transform 1 0 2512 0 1 1970
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1711653199
transform 1 0 2504 0 1 1970
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1711653199
transform 1 0 2496 0 1 1970
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1711653199
transform 1 0 2488 0 1 1970
box -8 -3 16 105
use FILL  FILL_1281
timestamp 1711653199
transform 1 0 2432 0 1 1970
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1711653199
transform 1 0 2424 0 1 1970
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1711653199
transform 1 0 2392 0 1 1970
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1711653199
transform 1 0 2336 0 1 1970
box -8 -3 16 105
use FILL  FILL_1285
timestamp 1711653199
transform 1 0 2328 0 1 1970
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1711653199
transform 1 0 2320 0 1 1970
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1711653199
transform 1 0 2296 0 1 1970
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1711653199
transform 1 0 2288 0 1 1970
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1711653199
transform 1 0 2256 0 1 1970
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1711653199
transform 1 0 2208 0 1 1970
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1711653199
transform 1 0 2200 0 1 1970
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1711653199
transform 1 0 2192 0 1 1970
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1711653199
transform 1 0 2152 0 1 1970
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1711653199
transform 1 0 2144 0 1 1970
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1711653199
transform 1 0 2080 0 1 1970
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1711653199
transform 1 0 2072 0 1 1970
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1711653199
transform 1 0 2064 0 1 1970
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1711653199
transform 1 0 2056 0 1 1970
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1711653199
transform 1 0 2000 0 1 1970
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1711653199
transform 1 0 1992 0 1 1970
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1711653199
transform 1 0 1960 0 1 1970
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1711653199
transform 1 0 1952 0 1 1970
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1711653199
transform 1 0 1912 0 1 1970
box -8 -3 16 105
use FILL  FILL_1304
timestamp 1711653199
transform 1 0 1904 0 1 1970
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1711653199
transform 1 0 1896 0 1 1970
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1711653199
transform 1 0 1888 0 1 1970
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1711653199
transform 1 0 1848 0 1 1970
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1711653199
transform 1 0 1840 0 1 1970
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1711653199
transform 1 0 1800 0 1 1970
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1711653199
transform 1 0 1792 0 1 1970
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1711653199
transform 1 0 1784 0 1 1970
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1711653199
transform 1 0 1720 0 1 1970
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1711653199
transform 1 0 1712 0 1 1970
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1711653199
transform 1 0 1688 0 1 1970
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1711653199
transform 1 0 1680 0 1 1970
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1711653199
transform 1 0 1672 0 1 1970
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1711653199
transform 1 0 1640 0 1 1970
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1711653199
transform 1 0 1632 0 1 1970
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1711653199
transform 1 0 1600 0 1 1970
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1711653199
transform 1 0 1592 0 1 1970
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1711653199
transform 1 0 1584 0 1 1970
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1711653199
transform 1 0 1576 0 1 1970
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1711653199
transform 1 0 1568 0 1 1970
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1711653199
transform 1 0 1520 0 1 1970
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1711653199
transform 1 0 1512 0 1 1970
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1711653199
transform 1 0 1504 0 1 1970
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1711653199
transform 1 0 1496 0 1 1970
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1711653199
transform 1 0 1488 0 1 1970
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1711653199
transform 1 0 1480 0 1 1970
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1711653199
transform 1 0 1440 0 1 1970
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1711653199
transform 1 0 1432 0 1 1970
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1711653199
transform 1 0 1424 0 1 1970
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1711653199
transform 1 0 1416 0 1 1970
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1711653199
transform 1 0 1408 0 1 1970
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1711653199
transform 1 0 1360 0 1 1970
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1711653199
transform 1 0 1352 0 1 1970
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1711653199
transform 1 0 1344 0 1 1970
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1711653199
transform 1 0 1336 0 1 1970
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1711653199
transform 1 0 1328 0 1 1970
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1711653199
transform 1 0 1320 0 1 1970
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1711653199
transform 1 0 1312 0 1 1970
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1711653199
transform 1 0 1256 0 1 1970
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1711653199
transform 1 0 1248 0 1 1970
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1711653199
transform 1 0 1200 0 1 1970
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1711653199
transform 1 0 1192 0 1 1970
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1711653199
transform 1 0 1184 0 1 1970
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1711653199
transform 1 0 1176 0 1 1970
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1711653199
transform 1 0 1168 0 1 1970
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1711653199
transform 1 0 1128 0 1 1970
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1711653199
transform 1 0 1120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1711653199
transform 1 0 1096 0 1 1970
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1711653199
transform 1 0 1088 0 1 1970
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1711653199
transform 1 0 1080 0 1 1970
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1711653199
transform 1 0 1056 0 1 1970
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1711653199
transform 1 0 1048 0 1 1970
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1711653199
transform 1 0 1040 0 1 1970
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1711653199
transform 1 0 1032 0 1 1970
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1711653199
transform 1 0 992 0 1 1970
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1711653199
transform 1 0 984 0 1 1970
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1711653199
transform 1 0 976 0 1 1970
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1711653199
transform 1 0 968 0 1 1970
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1711653199
transform 1 0 960 0 1 1970
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1711653199
transform 1 0 936 0 1 1970
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1711653199
transform 1 0 896 0 1 1970
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1711653199
transform 1 0 888 0 1 1970
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1711653199
transform 1 0 856 0 1 1970
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1711653199
transform 1 0 848 0 1 1970
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1711653199
transform 1 0 840 0 1 1970
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1711653199
transform 1 0 792 0 1 1970
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1711653199
transform 1 0 784 0 1 1970
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1711653199
transform 1 0 776 0 1 1970
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1711653199
transform 1 0 728 0 1 1970
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1711653199
transform 1 0 720 0 1 1970
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1711653199
transform 1 0 712 0 1 1970
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1711653199
transform 1 0 664 0 1 1970
box -8 -3 16 105
use FILL  FILL_1376
timestamp 1711653199
transform 1 0 656 0 1 1970
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1711653199
transform 1 0 648 0 1 1970
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1711653199
transform 1 0 608 0 1 1970
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1711653199
transform 1 0 600 0 1 1970
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1711653199
transform 1 0 592 0 1 1970
box -8 -3 16 105
use FILL  FILL_1381
timestamp 1711653199
transform 1 0 584 0 1 1970
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1711653199
transform 1 0 544 0 1 1970
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1711653199
transform 1 0 536 0 1 1970
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1711653199
transform 1 0 528 0 1 1970
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1711653199
transform 1 0 496 0 1 1970
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1711653199
transform 1 0 472 0 1 1970
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1711653199
transform 1 0 464 0 1 1970
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1711653199
transform 1 0 424 0 1 1970
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1711653199
transform 1 0 416 0 1 1970
box -8 -3 16 105
use FILL  FILL_1390
timestamp 1711653199
transform 1 0 384 0 1 1970
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1711653199
transform 1 0 376 0 1 1970
box -8 -3 16 105
use FILL  FILL_1392
timestamp 1711653199
transform 1 0 312 0 1 1970
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1711653199
transform 1 0 304 0 1 1970
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1711653199
transform 1 0 296 0 1 1970
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1711653199
transform 1 0 288 0 1 1970
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1711653199
transform 1 0 216 0 1 1970
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1711653199
transform 1 0 208 0 1 1970
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1711653199
transform 1 0 200 0 1 1970
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1711653199
transform 1 0 192 0 1 1970
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1711653199
transform 1 0 128 0 1 1970
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1711653199
transform 1 0 120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1711653199
transform 1 0 112 0 1 1970
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1711653199
transform 1 0 72 0 1 1970
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1711653199
transform 1 0 3128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1711653199
transform 1 0 3088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1711653199
transform 1 0 3080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1711653199
transform 1 0 3072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1711653199
transform 1 0 3024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1711653199
transform 1 0 2992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1711653199
transform 1 0 2984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1711653199
transform 1 0 2976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1711653199
transform 1 0 2912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1711653199
transform 1 0 2904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1711653199
transform 1 0 2896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1711653199
transform 1 0 2888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1711653199
transform 1 0 2816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1711653199
transform 1 0 2808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1711653199
transform 1 0 2800 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1711653199
transform 1 0 2792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1711653199
transform 1 0 2720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1711653199
transform 1 0 2712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1711653199
transform 1 0 2704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1711653199
transform 1 0 2672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1711653199
transform 1 0 2608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1711653199
transform 1 0 2600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1711653199
transform 1 0 2592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1711653199
transform 1 0 2552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1711653199
transform 1 0 2512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1711653199
transform 1 0 2488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1430
timestamp 1711653199
transform 1 0 2480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1711653199
transform 1 0 2432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1711653199
transform 1 0 2424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1711653199
transform 1 0 2416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1711653199
transform 1 0 2344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1711653199
transform 1 0 2336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1711653199
transform 1 0 2328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1711653199
transform 1 0 2264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1711653199
transform 1 0 2256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1711653199
transform 1 0 2184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1711653199
transform 1 0 2176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1711653199
transform 1 0 2168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1711653199
transform 1 0 2080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1711653199
transform 1 0 2072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1711653199
transform 1 0 2064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1711653199
transform 1 0 2056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1711653199
transform 1 0 1960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1711653199
transform 1 0 1952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1711653199
transform 1 0 1944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1711653199
transform 1 0 1936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1711653199
transform 1 0 1888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1711653199
transform 1 0 1848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1711653199
transform 1 0 1840 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1453
timestamp 1711653199
transform 1 0 1832 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1711653199
transform 1 0 1792 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1711653199
transform 1 0 1784 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1711653199
transform 1 0 1736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1711653199
transform 1 0 1648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1711653199
transform 1 0 1640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1711653199
transform 1 0 1632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1711653199
transform 1 0 1624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1711653199
transform 1 0 1584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1711653199
transform 1 0 1576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1711653199
transform 1 0 1544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1711653199
transform 1 0 1536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1711653199
transform 1 0 1528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1711653199
transform 1 0 1520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1711653199
transform 1 0 1512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1711653199
transform 1 0 1488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1711653199
transform 1 0 1448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1711653199
transform 1 0 1440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1711653199
transform 1 0 1432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1711653199
transform 1 0 1424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1711653199
transform 1 0 1416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1711653199
transform 1 0 1384 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1711653199
transform 1 0 1376 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1711653199
transform 1 0 1368 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1711653199
transform 1 0 1328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1711653199
transform 1 0 1320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1711653199
transform 1 0 1312 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1711653199
transform 1 0 1272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1711653199
transform 1 0 1264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1711653199
transform 1 0 1256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1711653199
transform 1 0 1184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1711653199
transform 1 0 1176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1711653199
transform 1 0 1168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1711653199
transform 1 0 1160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1711653199
transform 1 0 1120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1711653199
transform 1 0 1112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1711653199
transform 1 0 1104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1490
timestamp 1711653199
transform 1 0 1072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1711653199
transform 1 0 1064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1711653199
transform 1 0 1040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1711653199
transform 1 0 1032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1711653199
transform 1 0 1024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1711653199
transform 1 0 1016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1711653199
transform 1 0 1008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1711653199
transform 1 0 960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1711653199
transform 1 0 952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1711653199
transform 1 0 944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1711653199
transform 1 0 936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1711653199
transform 1 0 896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1711653199
transform 1 0 888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1711653199
transform 1 0 856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1711653199
transform 1 0 848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1711653199
transform 1 0 840 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1711653199
transform 1 0 816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1711653199
transform 1 0 808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1508
timestamp 1711653199
transform 1 0 768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1711653199
transform 1 0 760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1510
timestamp 1711653199
transform 1 0 752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1711653199
transform 1 0 744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1711653199
transform 1 0 704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1711653199
transform 1 0 696 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1514
timestamp 1711653199
transform 1 0 656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1711653199
transform 1 0 648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1711653199
transform 1 0 640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1711653199
transform 1 0 600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1711653199
transform 1 0 592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1711653199
transform 1 0 584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1520
timestamp 1711653199
transform 1 0 560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1711653199
transform 1 0 520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1711653199
transform 1 0 512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1711653199
transform 1 0 472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1711653199
transform 1 0 432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1711653199
transform 1 0 424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1711653199
transform 1 0 360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1711653199
transform 1 0 352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1711653199
transform 1 0 344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1711653199
transform 1 0 288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1711653199
transform 1 0 216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1711653199
transform 1 0 208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1711653199
transform 1 0 160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1711653199
transform 1 0 152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1711653199
transform 1 0 144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1711653199
transform 1 0 136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1711653199
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1711653199
transform 1 0 3392 0 1 1770
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1711653199
transform 1 0 3384 0 1 1770
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1711653199
transform 1 0 3376 0 1 1770
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1711653199
transform 1 0 3368 0 1 1770
box -8 -3 16 105
use FILL  FILL_1541
timestamp 1711653199
transform 1 0 3360 0 1 1770
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1711653199
transform 1 0 3336 0 1 1770
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1711653199
transform 1 0 3272 0 1 1770
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1711653199
transform 1 0 3264 0 1 1770
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1711653199
transform 1 0 3256 0 1 1770
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1711653199
transform 1 0 3248 0 1 1770
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1711653199
transform 1 0 3240 0 1 1770
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1711653199
transform 1 0 3176 0 1 1770
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1711653199
transform 1 0 3168 0 1 1770
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1711653199
transform 1 0 3144 0 1 1770
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1711653199
transform 1 0 3136 0 1 1770
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1711653199
transform 1 0 3128 0 1 1770
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1711653199
transform 1 0 3120 0 1 1770
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1711653199
transform 1 0 3112 0 1 1770
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1711653199
transform 1 0 3056 0 1 1770
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1711653199
transform 1 0 3048 0 1 1770
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1711653199
transform 1 0 3040 0 1 1770
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1711653199
transform 1 0 3032 0 1 1770
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1711653199
transform 1 0 3024 0 1 1770
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1711653199
transform 1 0 2960 0 1 1770
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1711653199
transform 1 0 2952 0 1 1770
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1711653199
transform 1 0 2944 0 1 1770
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1711653199
transform 1 0 2936 0 1 1770
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1711653199
transform 1 0 2896 0 1 1770
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1711653199
transform 1 0 2888 0 1 1770
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1711653199
transform 1 0 2880 0 1 1770
box -8 -3 16 105
use FILL  FILL_1567
timestamp 1711653199
transform 1 0 2824 0 1 1770
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1711653199
transform 1 0 2816 0 1 1770
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1711653199
transform 1 0 2808 0 1 1770
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1711653199
transform 1 0 2800 0 1 1770
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1711653199
transform 1 0 2728 0 1 1770
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1711653199
transform 1 0 2720 0 1 1770
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1711653199
transform 1 0 2712 0 1 1770
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1711653199
transform 1 0 2704 0 1 1770
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1711653199
transform 1 0 2696 0 1 1770
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1711653199
transform 1 0 2624 0 1 1770
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1711653199
transform 1 0 2616 0 1 1770
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1711653199
transform 1 0 2608 0 1 1770
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1711653199
transform 1 0 2600 0 1 1770
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1711653199
transform 1 0 2528 0 1 1770
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1711653199
transform 1 0 2520 0 1 1770
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1711653199
transform 1 0 2512 0 1 1770
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1711653199
transform 1 0 2504 0 1 1770
box -8 -3 16 105
use FILL  FILL_1584
timestamp 1711653199
transform 1 0 2496 0 1 1770
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1711653199
transform 1 0 2488 0 1 1770
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1711653199
transform 1 0 2416 0 1 1770
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1711653199
transform 1 0 2408 0 1 1770
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1711653199
transform 1 0 2400 0 1 1770
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1711653199
transform 1 0 2392 0 1 1770
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1711653199
transform 1 0 2320 0 1 1770
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1711653199
transform 1 0 2312 0 1 1770
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1711653199
transform 1 0 2304 0 1 1770
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1711653199
transform 1 0 2296 0 1 1770
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1711653199
transform 1 0 2288 0 1 1770
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1711653199
transform 1 0 2216 0 1 1770
box -8 -3 16 105
use FILL  FILL_1596
timestamp 1711653199
transform 1 0 2208 0 1 1770
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1711653199
transform 1 0 2200 0 1 1770
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1711653199
transform 1 0 2192 0 1 1770
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1711653199
transform 1 0 2152 0 1 1770
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1711653199
transform 1 0 2112 0 1 1770
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1711653199
transform 1 0 2104 0 1 1770
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1711653199
transform 1 0 2096 0 1 1770
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1711653199
transform 1 0 2072 0 1 1770
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1711653199
transform 1 0 2064 0 1 1770
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1711653199
transform 1 0 2056 0 1 1770
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1711653199
transform 1 0 2000 0 1 1770
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1711653199
transform 1 0 1992 0 1 1770
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1711653199
transform 1 0 1984 0 1 1770
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1711653199
transform 1 0 1976 0 1 1770
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1711653199
transform 1 0 1952 0 1 1770
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1711653199
transform 1 0 1944 0 1 1770
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1711653199
transform 1 0 1904 0 1 1770
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1711653199
transform 1 0 1896 0 1 1770
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1711653199
transform 1 0 1888 0 1 1770
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1711653199
transform 1 0 1880 0 1 1770
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1711653199
transform 1 0 1872 0 1 1770
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1711653199
transform 1 0 1864 0 1 1770
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1711653199
transform 1 0 1816 0 1 1770
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1711653199
transform 1 0 1808 0 1 1770
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1711653199
transform 1 0 1800 0 1 1770
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1711653199
transform 1 0 1792 0 1 1770
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1711653199
transform 1 0 1784 0 1 1770
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1711653199
transform 1 0 1776 0 1 1770
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1711653199
transform 1 0 1768 0 1 1770
box -8 -3 16 105
use FILL  FILL_1625
timestamp 1711653199
transform 1 0 1720 0 1 1770
box -8 -3 16 105
use FILL  FILL_1626
timestamp 1711653199
transform 1 0 1712 0 1 1770
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1711653199
transform 1 0 1704 0 1 1770
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1711653199
transform 1 0 1696 0 1 1770
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1711653199
transform 1 0 1664 0 1 1770
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1711653199
transform 1 0 1656 0 1 1770
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1711653199
transform 1 0 1648 0 1 1770
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1711653199
transform 1 0 1616 0 1 1770
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1711653199
transform 1 0 1608 0 1 1770
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1711653199
transform 1 0 1600 0 1 1770
box -8 -3 16 105
use FILL  FILL_1635
timestamp 1711653199
transform 1 0 1592 0 1 1770
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1711653199
transform 1 0 1584 0 1 1770
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1711653199
transform 1 0 1576 0 1 1770
box -8 -3 16 105
use FILL  FILL_1638
timestamp 1711653199
transform 1 0 1536 0 1 1770
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1711653199
transform 1 0 1528 0 1 1770
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1711653199
transform 1 0 1520 0 1 1770
box -8 -3 16 105
use FILL  FILL_1641
timestamp 1711653199
transform 1 0 1512 0 1 1770
box -8 -3 16 105
use FILL  FILL_1642
timestamp 1711653199
transform 1 0 1480 0 1 1770
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1711653199
transform 1 0 1472 0 1 1770
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1711653199
transform 1 0 1464 0 1 1770
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1711653199
transform 1 0 1456 0 1 1770
box -8 -3 16 105
use FILL  FILL_1646
timestamp 1711653199
transform 1 0 1448 0 1 1770
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1711653199
transform 1 0 1408 0 1 1770
box -8 -3 16 105
use FILL  FILL_1648
timestamp 1711653199
transform 1 0 1400 0 1 1770
box -8 -3 16 105
use FILL  FILL_1649
timestamp 1711653199
transform 1 0 1392 0 1 1770
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1711653199
transform 1 0 1384 0 1 1770
box -8 -3 16 105
use FILL  FILL_1651
timestamp 1711653199
transform 1 0 1376 0 1 1770
box -8 -3 16 105
use FILL  FILL_1652
timestamp 1711653199
transform 1 0 1336 0 1 1770
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1711653199
transform 1 0 1328 0 1 1770
box -8 -3 16 105
use FILL  FILL_1654
timestamp 1711653199
transform 1 0 1320 0 1 1770
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1711653199
transform 1 0 1312 0 1 1770
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1711653199
transform 1 0 1304 0 1 1770
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1711653199
transform 1 0 1264 0 1 1770
box -8 -3 16 105
use FILL  FILL_1658
timestamp 1711653199
transform 1 0 1256 0 1 1770
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1711653199
transform 1 0 1248 0 1 1770
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1711653199
transform 1 0 1240 0 1 1770
box -8 -3 16 105
use FILL  FILL_1661
timestamp 1711653199
transform 1 0 1232 0 1 1770
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1711653199
transform 1 0 1192 0 1 1770
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1711653199
transform 1 0 1184 0 1 1770
box -8 -3 16 105
use FILL  FILL_1664
timestamp 1711653199
transform 1 0 1144 0 1 1770
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1711653199
transform 1 0 1136 0 1 1770
box -8 -3 16 105
use FILL  FILL_1666
timestamp 1711653199
transform 1 0 1128 0 1 1770
box -8 -3 16 105
use FILL  FILL_1667
timestamp 1711653199
transform 1 0 1120 0 1 1770
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1711653199
transform 1 0 1112 0 1 1770
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1711653199
transform 1 0 1072 0 1 1770
box -8 -3 16 105
use FILL  FILL_1670
timestamp 1711653199
transform 1 0 1064 0 1 1770
box -8 -3 16 105
use FILL  FILL_1671
timestamp 1711653199
transform 1 0 1056 0 1 1770
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1711653199
transform 1 0 1048 0 1 1770
box -8 -3 16 105
use FILL  FILL_1673
timestamp 1711653199
transform 1 0 1040 0 1 1770
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1711653199
transform 1 0 1000 0 1 1770
box -8 -3 16 105
use FILL  FILL_1675
timestamp 1711653199
transform 1 0 992 0 1 1770
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1711653199
transform 1 0 984 0 1 1770
box -8 -3 16 105
use FILL  FILL_1677
timestamp 1711653199
transform 1 0 976 0 1 1770
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1711653199
transform 1 0 968 0 1 1770
box -8 -3 16 105
use FILL  FILL_1679
timestamp 1711653199
transform 1 0 960 0 1 1770
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1711653199
transform 1 0 920 0 1 1770
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1711653199
transform 1 0 888 0 1 1770
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1711653199
transform 1 0 880 0 1 1770
box -8 -3 16 105
use FILL  FILL_1683
timestamp 1711653199
transform 1 0 872 0 1 1770
box -8 -3 16 105
use FILL  FILL_1684
timestamp 1711653199
transform 1 0 840 0 1 1770
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1711653199
transform 1 0 832 0 1 1770
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1711653199
transform 1 0 824 0 1 1770
box -8 -3 16 105
use FILL  FILL_1687
timestamp 1711653199
transform 1 0 784 0 1 1770
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1711653199
transform 1 0 776 0 1 1770
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1711653199
transform 1 0 768 0 1 1770
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1711653199
transform 1 0 760 0 1 1770
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1711653199
transform 1 0 720 0 1 1770
box -8 -3 16 105
use FILL  FILL_1692
timestamp 1711653199
transform 1 0 712 0 1 1770
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1711653199
transform 1 0 704 0 1 1770
box -8 -3 16 105
use FILL  FILL_1694
timestamp 1711653199
transform 1 0 696 0 1 1770
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1711653199
transform 1 0 688 0 1 1770
box -8 -3 16 105
use FILL  FILL_1696
timestamp 1711653199
transform 1 0 648 0 1 1770
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1711653199
transform 1 0 640 0 1 1770
box -8 -3 16 105
use FILL  FILL_1698
timestamp 1711653199
transform 1 0 632 0 1 1770
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1711653199
transform 1 0 592 0 1 1770
box -8 -3 16 105
use FILL  FILL_1700
timestamp 1711653199
transform 1 0 584 0 1 1770
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1711653199
transform 1 0 576 0 1 1770
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1711653199
transform 1 0 536 0 1 1770
box -8 -3 16 105
use FILL  FILL_1703
timestamp 1711653199
transform 1 0 504 0 1 1770
box -8 -3 16 105
use FILL  FILL_1704
timestamp 1711653199
transform 1 0 496 0 1 1770
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1711653199
transform 1 0 464 0 1 1770
box -8 -3 16 105
use FILL  FILL_1706
timestamp 1711653199
transform 1 0 456 0 1 1770
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1711653199
transform 1 0 448 0 1 1770
box -8 -3 16 105
use FILL  FILL_1708
timestamp 1711653199
transform 1 0 376 0 1 1770
box -8 -3 16 105
use FILL  FILL_1709
timestamp 1711653199
transform 1 0 368 0 1 1770
box -8 -3 16 105
use FILL  FILL_1710
timestamp 1711653199
transform 1 0 360 0 1 1770
box -8 -3 16 105
use FILL  FILL_1711
timestamp 1711653199
transform 1 0 296 0 1 1770
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1711653199
transform 1 0 288 0 1 1770
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1711653199
transform 1 0 280 0 1 1770
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1711653199
transform 1 0 208 0 1 1770
box -8 -3 16 105
use FILL  FILL_1715
timestamp 1711653199
transform 1 0 200 0 1 1770
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1711653199
transform 1 0 160 0 1 1770
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1711653199
transform 1 0 152 0 1 1770
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1711653199
transform 1 0 144 0 1 1770
box -8 -3 16 105
use FILL  FILL_1719
timestamp 1711653199
transform 1 0 136 0 1 1770
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1711653199
transform 1 0 80 0 1 1770
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1711653199
transform 1 0 72 0 1 1770
box -8 -3 16 105
use FILL  FILL_1722
timestamp 1711653199
transform 1 0 3392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1711653199
transform 1 0 3384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1711653199
transform 1 0 3344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1725
timestamp 1711653199
transform 1 0 3336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1711653199
transform 1 0 3328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1711653199
transform 1 0 3288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1711653199
transform 1 0 3280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1729
timestamp 1711653199
transform 1 0 3272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1711653199
transform 1 0 3216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1711653199
transform 1 0 3208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1711653199
transform 1 0 3200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1711653199
transform 1 0 3192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1734
timestamp 1711653199
transform 1 0 3128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1711653199
transform 1 0 3120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1736
timestamp 1711653199
transform 1 0 3112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1737
timestamp 1711653199
transform 1 0 3104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1711653199
transform 1 0 3064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1711653199
transform 1 0 3056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1740
timestamp 1711653199
transform 1 0 3016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1711653199
transform 1 0 3008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1742
timestamp 1711653199
transform 1 0 3000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1711653199
transform 1 0 2992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1711653199
transform 1 0 2944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1745
timestamp 1711653199
transform 1 0 2936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1746
timestamp 1711653199
transform 1 0 2928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1711653199
transform 1 0 2904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1711653199
transform 1 0 2896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1749
timestamp 1711653199
transform 1 0 2848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1711653199
transform 1 0 2840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1751
timestamp 1711653199
transform 1 0 2832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1711653199
transform 1 0 2824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1753
timestamp 1711653199
transform 1 0 2816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1711653199
transform 1 0 2768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1755
timestamp 1711653199
transform 1 0 2728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1711653199
transform 1 0 2720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1757
timestamp 1711653199
transform 1 0 2712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1711653199
transform 1 0 2704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1711653199
transform 1 0 2696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1760
timestamp 1711653199
transform 1 0 2664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1761
timestamp 1711653199
transform 1 0 2624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1762
timestamp 1711653199
transform 1 0 2616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1711653199
transform 1 0 2608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1764
timestamp 1711653199
transform 1 0 2600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1765
timestamp 1711653199
transform 1 0 2552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1711653199
transform 1 0 2544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1767
timestamp 1711653199
transform 1 0 2504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1711653199
transform 1 0 2496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1711653199
transform 1 0 2488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1770
timestamp 1711653199
transform 1 0 2480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1771
timestamp 1711653199
transform 1 0 2416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1772
timestamp 1711653199
transform 1 0 2408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1711653199
transform 1 0 2400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1774
timestamp 1711653199
transform 1 0 2392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1711653199
transform 1 0 2320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1776
timestamp 1711653199
transform 1 0 2312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1777
timestamp 1711653199
transform 1 0 2304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1711653199
transform 1 0 2296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1779
timestamp 1711653199
transform 1 0 2256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1711653199
transform 1 0 2216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1711653199
transform 1 0 2208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1711653199
transform 1 0 2184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1711653199
transform 1 0 2176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1784
timestamp 1711653199
transform 1 0 2168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1711653199
transform 1 0 2160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1786
timestamp 1711653199
transform 1 0 2096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1711653199
transform 1 0 2088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1788
timestamp 1711653199
transform 1 0 2080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1789
timestamp 1711653199
transform 1 0 2008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1790
timestamp 1711653199
transform 1 0 2000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1711653199
transform 1 0 1992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1792
timestamp 1711653199
transform 1 0 1952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1793
timestamp 1711653199
transform 1 0 1944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1711653199
transform 1 0 1904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1795
timestamp 1711653199
transform 1 0 1896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1711653199
transform 1 0 1888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1711653199
transform 1 0 1848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1711653199
transform 1 0 1840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1799
timestamp 1711653199
transform 1 0 1832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1711653199
transform 1 0 1792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1711653199
transform 1 0 1784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1711653199
transform 1 0 1776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1711653199
transform 1 0 1768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1711653199
transform 1 0 1760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1711653199
transform 1 0 1720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1711653199
transform 1 0 1712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1807
timestamp 1711653199
transform 1 0 1704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1711653199
transform 1 0 1696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1809
timestamp 1711653199
transform 1 0 1688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1711653199
transform 1 0 1680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1711653199
transform 1 0 1648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1812
timestamp 1711653199
transform 1 0 1640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1711653199
transform 1 0 1632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1711653199
transform 1 0 1624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1711653199
transform 1 0 1584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1711653199
transform 1 0 1576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1817
timestamp 1711653199
transform 1 0 1568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1818
timestamp 1711653199
transform 1 0 1560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1711653199
transform 1 0 1552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1820
timestamp 1711653199
transform 1 0 1544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1711653199
transform 1 0 1520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1711653199
transform 1 0 1512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1823
timestamp 1711653199
transform 1 0 1488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1824
timestamp 1711653199
transform 1 0 1480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1825
timestamp 1711653199
transform 1 0 1472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1711653199
transform 1 0 1464 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1827
timestamp 1711653199
transform 1 0 1456 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1711653199
transform 1 0 1424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1829
timestamp 1711653199
transform 1 0 1416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1830
timestamp 1711653199
transform 1 0 1408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1711653199
transform 1 0 1400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1711653199
transform 1 0 1360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1711653199
transform 1 0 1352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1711653199
transform 1 0 1344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1835
timestamp 1711653199
transform 1 0 1336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1711653199
transform 1 0 1328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1837
timestamp 1711653199
transform 1 0 1320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1711653199
transform 1 0 1312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1839
timestamp 1711653199
transform 1 0 1272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1711653199
transform 1 0 1264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1711653199
transform 1 0 1256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1711653199
transform 1 0 1248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1711653199
transform 1 0 1240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1711653199
transform 1 0 1232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1711653199
transform 1 0 1224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1711653199
transform 1 0 1184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1711653199
transform 1 0 1176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1848
timestamp 1711653199
transform 1 0 1168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1711653199
transform 1 0 1160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1711653199
transform 1 0 1152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1711653199
transform 1 0 1112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1711653199
transform 1 0 1104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1711653199
transform 1 0 1096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1854
timestamp 1711653199
transform 1 0 1088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1855
timestamp 1711653199
transform 1 0 1080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1711653199
transform 1 0 1072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1857
timestamp 1711653199
transform 1 0 1064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1711653199
transform 1 0 1056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1711653199
transform 1 0 1016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1860
timestamp 1711653199
transform 1 0 1008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1711653199
transform 1 0 1000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1711653199
transform 1 0 992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1863
timestamp 1711653199
transform 1 0 984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1711653199
transform 1 0 976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1711653199
transform 1 0 936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1711653199
transform 1 0 928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1711653199
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1711653199
transform 1 0 912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1869
timestamp 1711653199
transform 1 0 904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1870
timestamp 1711653199
transform 1 0 896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1871
timestamp 1711653199
transform 1 0 864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1711653199
transform 1 0 856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1873
timestamp 1711653199
transform 1 0 848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1874
timestamp 1711653199
transform 1 0 840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1711653199
transform 1 0 800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1711653199
transform 1 0 792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1877
timestamp 1711653199
transform 1 0 784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1711653199
transform 1 0 776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1711653199
transform 1 0 768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1711653199
transform 1 0 760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1711653199
transform 1 0 728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1882
timestamp 1711653199
transform 1 0 720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1711653199
transform 1 0 712 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1884
timestamp 1711653199
transform 1 0 704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1885
timestamp 1711653199
transform 1 0 664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1886
timestamp 1711653199
transform 1 0 656 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1711653199
transform 1 0 624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1888
timestamp 1711653199
transform 1 0 616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1889
timestamp 1711653199
transform 1 0 608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1711653199
transform 1 0 600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1891
timestamp 1711653199
transform 1 0 592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1711653199
transform 1 0 520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1893
timestamp 1711653199
transform 1 0 512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1894
timestamp 1711653199
transform 1 0 504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1895
timestamp 1711653199
transform 1 0 496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1711653199
transform 1 0 488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1711653199
transform 1 0 480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1898
timestamp 1711653199
transform 1 0 392 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1711653199
transform 1 0 384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1900
timestamp 1711653199
transform 1 0 376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1711653199
transform 1 0 368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1711653199
transform 1 0 360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1711653199
transform 1 0 288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1904
timestamp 1711653199
transform 1 0 280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1711653199
transform 1 0 272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1711653199
transform 1 0 264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1907
timestamp 1711653199
transform 1 0 200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1908
timestamp 1711653199
transform 1 0 152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1909
timestamp 1711653199
transform 1 0 144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1711653199
transform 1 0 136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1911
timestamp 1711653199
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1711653199
transform 1 0 3392 0 1 1570
box -8 -3 16 105
use FILL  FILL_1913
timestamp 1711653199
transform 1 0 3384 0 1 1570
box -8 -3 16 105
use FILL  FILL_1914
timestamp 1711653199
transform 1 0 3376 0 1 1570
box -8 -3 16 105
use FILL  FILL_1915
timestamp 1711653199
transform 1 0 3368 0 1 1570
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1711653199
transform 1 0 3304 0 1 1570
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1711653199
transform 1 0 3296 0 1 1570
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1711653199
transform 1 0 3288 0 1 1570
box -8 -3 16 105
use FILL  FILL_1919
timestamp 1711653199
transform 1 0 3280 0 1 1570
box -8 -3 16 105
use FILL  FILL_1920
timestamp 1711653199
transform 1 0 3272 0 1 1570
box -8 -3 16 105
use FILL  FILL_1921
timestamp 1711653199
transform 1 0 3208 0 1 1570
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1711653199
transform 1 0 3200 0 1 1570
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1711653199
transform 1 0 3192 0 1 1570
box -8 -3 16 105
use FILL  FILL_1924
timestamp 1711653199
transform 1 0 3184 0 1 1570
box -8 -3 16 105
use FILL  FILL_1925
timestamp 1711653199
transform 1 0 3176 0 1 1570
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1711653199
transform 1 0 3120 0 1 1570
box -8 -3 16 105
use FILL  FILL_1927
timestamp 1711653199
transform 1 0 3088 0 1 1570
box -8 -3 16 105
use FILL  FILL_1928
timestamp 1711653199
transform 1 0 3080 0 1 1570
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1711653199
transform 1 0 3072 0 1 1570
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1711653199
transform 1 0 3016 0 1 1570
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1711653199
transform 1 0 3008 0 1 1570
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1711653199
transform 1 0 2984 0 1 1570
box -8 -3 16 105
use FILL  FILL_1933
timestamp 1711653199
transform 1 0 2976 0 1 1570
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1711653199
transform 1 0 2968 0 1 1570
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1711653199
transform 1 0 2960 0 1 1570
box -8 -3 16 105
use FILL  FILL_1936
timestamp 1711653199
transform 1 0 2920 0 1 1570
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1711653199
transform 1 0 2880 0 1 1570
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1711653199
transform 1 0 2872 0 1 1570
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1711653199
transform 1 0 2864 0 1 1570
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1711653199
transform 1 0 2856 0 1 1570
box -8 -3 16 105
use FILL  FILL_1941
timestamp 1711653199
transform 1 0 2816 0 1 1570
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1711653199
transform 1 0 2768 0 1 1570
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1711653199
transform 1 0 2760 0 1 1570
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1711653199
transform 1 0 2752 0 1 1570
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1711653199
transform 1 0 2744 0 1 1570
box -8 -3 16 105
use FILL  FILL_1946
timestamp 1711653199
transform 1 0 2736 0 1 1570
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1711653199
transform 1 0 2664 0 1 1570
box -8 -3 16 105
use FILL  FILL_1948
timestamp 1711653199
transform 1 0 2656 0 1 1570
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1711653199
transform 1 0 2648 0 1 1570
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1711653199
transform 1 0 2640 0 1 1570
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1711653199
transform 1 0 2592 0 1 1570
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1711653199
transform 1 0 2584 0 1 1570
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1711653199
transform 1 0 2536 0 1 1570
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1711653199
transform 1 0 2528 0 1 1570
box -8 -3 16 105
use FILL  FILL_1955
timestamp 1711653199
transform 1 0 2520 0 1 1570
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1711653199
transform 1 0 2512 0 1 1570
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1711653199
transform 1 0 2472 0 1 1570
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1711653199
transform 1 0 2464 0 1 1570
box -8 -3 16 105
use FILL  FILL_1959
timestamp 1711653199
transform 1 0 2424 0 1 1570
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1711653199
transform 1 0 2416 0 1 1570
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1711653199
transform 1 0 2408 0 1 1570
box -8 -3 16 105
use FILL  FILL_1962
timestamp 1711653199
transform 1 0 2400 0 1 1570
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1711653199
transform 1 0 2360 0 1 1570
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1711653199
transform 1 0 2352 0 1 1570
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1711653199
transform 1 0 2344 0 1 1570
box -8 -3 16 105
use FILL  FILL_1966
timestamp 1711653199
transform 1 0 2296 0 1 1570
box -8 -3 16 105
use FILL  FILL_1967
timestamp 1711653199
transform 1 0 2288 0 1 1570
box -8 -3 16 105
use FILL  FILL_1968
timestamp 1711653199
transform 1 0 2240 0 1 1570
box -8 -3 16 105
use FILL  FILL_1969
timestamp 1711653199
transform 1 0 2232 0 1 1570
box -8 -3 16 105
use FILL  FILL_1970
timestamp 1711653199
transform 1 0 2200 0 1 1570
box -8 -3 16 105
use FILL  FILL_1971
timestamp 1711653199
transform 1 0 2168 0 1 1570
box -8 -3 16 105
use FILL  FILL_1972
timestamp 1711653199
transform 1 0 2160 0 1 1570
box -8 -3 16 105
use FILL  FILL_1973
timestamp 1711653199
transform 1 0 2120 0 1 1570
box -8 -3 16 105
use FILL  FILL_1974
timestamp 1711653199
transform 1 0 2072 0 1 1570
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1711653199
transform 1 0 2064 0 1 1570
box -8 -3 16 105
use FILL  FILL_1976
timestamp 1711653199
transform 1 0 2056 0 1 1570
box -8 -3 16 105
use FILL  FILL_1977
timestamp 1711653199
transform 1 0 2016 0 1 1570
box -8 -3 16 105
use FILL  FILL_1978
timestamp 1711653199
transform 1 0 1984 0 1 1570
box -8 -3 16 105
use FILL  FILL_1979
timestamp 1711653199
transform 1 0 1944 0 1 1570
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1711653199
transform 1 0 1936 0 1 1570
box -8 -3 16 105
use FILL  FILL_1981
timestamp 1711653199
transform 1 0 1928 0 1 1570
box -8 -3 16 105
use FILL  FILL_1982
timestamp 1711653199
transform 1 0 1896 0 1 1570
box -8 -3 16 105
use FILL  FILL_1983
timestamp 1711653199
transform 1 0 1888 0 1 1570
box -8 -3 16 105
use FILL  FILL_1984
timestamp 1711653199
transform 1 0 1840 0 1 1570
box -8 -3 16 105
use FILL  FILL_1985
timestamp 1711653199
transform 1 0 1832 0 1 1570
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1711653199
transform 1 0 1824 0 1 1570
box -8 -3 16 105
use FILL  FILL_1987
timestamp 1711653199
transform 1 0 1816 0 1 1570
box -8 -3 16 105
use FILL  FILL_1988
timestamp 1711653199
transform 1 0 1808 0 1 1570
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1711653199
transform 1 0 1800 0 1 1570
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1711653199
transform 1 0 1760 0 1 1570
box -8 -3 16 105
use FILL  FILL_1991
timestamp 1711653199
transform 1 0 1752 0 1 1570
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1711653199
transform 1 0 1720 0 1 1570
box -8 -3 16 105
use FILL  FILL_1993
timestamp 1711653199
transform 1 0 1712 0 1 1570
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1711653199
transform 1 0 1704 0 1 1570
box -8 -3 16 105
use FILL  FILL_1995
timestamp 1711653199
transform 1 0 1696 0 1 1570
box -8 -3 16 105
use FILL  FILL_1996
timestamp 1711653199
transform 1 0 1648 0 1 1570
box -8 -3 16 105
use FILL  FILL_1997
timestamp 1711653199
transform 1 0 1640 0 1 1570
box -8 -3 16 105
use FILL  FILL_1998
timestamp 1711653199
transform 1 0 1632 0 1 1570
box -8 -3 16 105
use FILL  FILL_1999
timestamp 1711653199
transform 1 0 1624 0 1 1570
box -8 -3 16 105
use FILL  FILL_2000
timestamp 1711653199
transform 1 0 1584 0 1 1570
box -8 -3 16 105
use FILL  FILL_2001
timestamp 1711653199
transform 1 0 1576 0 1 1570
box -8 -3 16 105
use FILL  FILL_2002
timestamp 1711653199
transform 1 0 1568 0 1 1570
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1711653199
transform 1 0 1528 0 1 1570
box -8 -3 16 105
use FILL  FILL_2004
timestamp 1711653199
transform 1 0 1520 0 1 1570
box -8 -3 16 105
use FILL  FILL_2005
timestamp 1711653199
transform 1 0 1512 0 1 1570
box -8 -3 16 105
use FILL  FILL_2006
timestamp 1711653199
transform 1 0 1504 0 1 1570
box -8 -3 16 105
use FILL  FILL_2007
timestamp 1711653199
transform 1 0 1464 0 1 1570
box -8 -3 16 105
use FILL  FILL_2008
timestamp 1711653199
transform 1 0 1456 0 1 1570
box -8 -3 16 105
use FILL  FILL_2009
timestamp 1711653199
transform 1 0 1448 0 1 1570
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1711653199
transform 1 0 1440 0 1 1570
box -8 -3 16 105
use FILL  FILL_2011
timestamp 1711653199
transform 1 0 1432 0 1 1570
box -8 -3 16 105
use FILL  FILL_2012
timestamp 1711653199
transform 1 0 1384 0 1 1570
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1711653199
transform 1 0 1376 0 1 1570
box -8 -3 16 105
use FILL  FILL_2014
timestamp 1711653199
transform 1 0 1368 0 1 1570
box -8 -3 16 105
use FILL  FILL_2015
timestamp 1711653199
transform 1 0 1360 0 1 1570
box -8 -3 16 105
use FILL  FILL_2016
timestamp 1711653199
transform 1 0 1352 0 1 1570
box -8 -3 16 105
use FILL  FILL_2017
timestamp 1711653199
transform 1 0 1312 0 1 1570
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1711653199
transform 1 0 1304 0 1 1570
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1711653199
transform 1 0 1296 0 1 1570
box -8 -3 16 105
use FILL  FILL_2020
timestamp 1711653199
transform 1 0 1288 0 1 1570
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1711653199
transform 1 0 1280 0 1 1570
box -8 -3 16 105
use FILL  FILL_2022
timestamp 1711653199
transform 1 0 1272 0 1 1570
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1711653199
transform 1 0 1264 0 1 1570
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1711653199
transform 1 0 1216 0 1 1570
box -8 -3 16 105
use FILL  FILL_2025
timestamp 1711653199
transform 1 0 1208 0 1 1570
box -8 -3 16 105
use FILL  FILL_2026
timestamp 1711653199
transform 1 0 1200 0 1 1570
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1711653199
transform 1 0 1192 0 1 1570
box -8 -3 16 105
use FILL  FILL_2028
timestamp 1711653199
transform 1 0 1184 0 1 1570
box -8 -3 16 105
use FILL  FILL_2029
timestamp 1711653199
transform 1 0 1144 0 1 1570
box -8 -3 16 105
use FILL  FILL_2030
timestamp 1711653199
transform 1 0 1136 0 1 1570
box -8 -3 16 105
use FILL  FILL_2031
timestamp 1711653199
transform 1 0 1128 0 1 1570
box -8 -3 16 105
use FILL  FILL_2032
timestamp 1711653199
transform 1 0 1120 0 1 1570
box -8 -3 16 105
use FILL  FILL_2033
timestamp 1711653199
transform 1 0 1112 0 1 1570
box -8 -3 16 105
use FILL  FILL_2034
timestamp 1711653199
transform 1 0 1080 0 1 1570
box -8 -3 16 105
use FILL  FILL_2035
timestamp 1711653199
transform 1 0 1072 0 1 1570
box -8 -3 16 105
use FILL  FILL_2036
timestamp 1711653199
transform 1 0 1064 0 1 1570
box -8 -3 16 105
use FILL  FILL_2037
timestamp 1711653199
transform 1 0 1056 0 1 1570
box -8 -3 16 105
use FILL  FILL_2038
timestamp 1711653199
transform 1 0 1016 0 1 1570
box -8 -3 16 105
use FILL  FILL_2039
timestamp 1711653199
transform 1 0 1008 0 1 1570
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1711653199
transform 1 0 1000 0 1 1570
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1711653199
transform 1 0 992 0 1 1570
box -8 -3 16 105
use FILL  FILL_2042
timestamp 1711653199
transform 1 0 984 0 1 1570
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1711653199
transform 1 0 976 0 1 1570
box -8 -3 16 105
use FILL  FILL_2044
timestamp 1711653199
transform 1 0 928 0 1 1570
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1711653199
transform 1 0 920 0 1 1570
box -8 -3 16 105
use FILL  FILL_2046
timestamp 1711653199
transform 1 0 912 0 1 1570
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1711653199
transform 1 0 904 0 1 1570
box -8 -3 16 105
use FILL  FILL_2048
timestamp 1711653199
transform 1 0 896 0 1 1570
box -8 -3 16 105
use FILL  FILL_2049
timestamp 1711653199
transform 1 0 872 0 1 1570
box -8 -3 16 105
use FILL  FILL_2050
timestamp 1711653199
transform 1 0 864 0 1 1570
box -8 -3 16 105
use FILL  FILL_2051
timestamp 1711653199
transform 1 0 856 0 1 1570
box -8 -3 16 105
use FILL  FILL_2052
timestamp 1711653199
transform 1 0 816 0 1 1570
box -8 -3 16 105
use FILL  FILL_2053
timestamp 1711653199
transform 1 0 808 0 1 1570
box -8 -3 16 105
use FILL  FILL_2054
timestamp 1711653199
transform 1 0 800 0 1 1570
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1711653199
transform 1 0 792 0 1 1570
box -8 -3 16 105
use FILL  FILL_2056
timestamp 1711653199
transform 1 0 784 0 1 1570
box -8 -3 16 105
use FILL  FILL_2057
timestamp 1711653199
transform 1 0 744 0 1 1570
box -8 -3 16 105
use FILL  FILL_2058
timestamp 1711653199
transform 1 0 736 0 1 1570
box -8 -3 16 105
use FILL  FILL_2059
timestamp 1711653199
transform 1 0 728 0 1 1570
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1711653199
transform 1 0 720 0 1 1570
box -8 -3 16 105
use FILL  FILL_2061
timestamp 1711653199
transform 1 0 712 0 1 1570
box -8 -3 16 105
use FILL  FILL_2062
timestamp 1711653199
transform 1 0 672 0 1 1570
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1711653199
transform 1 0 632 0 1 1570
box -8 -3 16 105
use FILL  FILL_2064
timestamp 1711653199
transform 1 0 624 0 1 1570
box -8 -3 16 105
use FILL  FILL_2065
timestamp 1711653199
transform 1 0 616 0 1 1570
box -8 -3 16 105
use FILL  FILL_2066
timestamp 1711653199
transform 1 0 576 0 1 1570
box -8 -3 16 105
use FILL  FILL_2067
timestamp 1711653199
transform 1 0 568 0 1 1570
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1711653199
transform 1 0 560 0 1 1570
box -8 -3 16 105
use FILL  FILL_2069
timestamp 1711653199
transform 1 0 512 0 1 1570
box -8 -3 16 105
use FILL  FILL_2070
timestamp 1711653199
transform 1 0 504 0 1 1570
box -8 -3 16 105
use FILL  FILL_2071
timestamp 1711653199
transform 1 0 496 0 1 1570
box -8 -3 16 105
use FILL  FILL_2072
timestamp 1711653199
transform 1 0 488 0 1 1570
box -8 -3 16 105
use FILL  FILL_2073
timestamp 1711653199
transform 1 0 448 0 1 1570
box -8 -3 16 105
use FILL  FILL_2074
timestamp 1711653199
transform 1 0 440 0 1 1570
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1711653199
transform 1 0 432 0 1 1570
box -8 -3 16 105
use FILL  FILL_2076
timestamp 1711653199
transform 1 0 400 0 1 1570
box -8 -3 16 105
use FILL  FILL_2077
timestamp 1711653199
transform 1 0 392 0 1 1570
box -8 -3 16 105
use FILL  FILL_2078
timestamp 1711653199
transform 1 0 384 0 1 1570
box -8 -3 16 105
use FILL  FILL_2079
timestamp 1711653199
transform 1 0 336 0 1 1570
box -8 -3 16 105
use FILL  FILL_2080
timestamp 1711653199
transform 1 0 328 0 1 1570
box -8 -3 16 105
use FILL  FILL_2081
timestamp 1711653199
transform 1 0 280 0 1 1570
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1711653199
transform 1 0 272 0 1 1570
box -8 -3 16 105
use FILL  FILL_2083
timestamp 1711653199
transform 1 0 264 0 1 1570
box -8 -3 16 105
use FILL  FILL_2084
timestamp 1711653199
transform 1 0 256 0 1 1570
box -8 -3 16 105
use FILL  FILL_2085
timestamp 1711653199
transform 1 0 224 0 1 1570
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1711653199
transform 1 0 176 0 1 1570
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1711653199
transform 1 0 168 0 1 1570
box -8 -3 16 105
use FILL  FILL_2088
timestamp 1711653199
transform 1 0 160 0 1 1570
box -8 -3 16 105
use FILL  FILL_2089
timestamp 1711653199
transform 1 0 152 0 1 1570
box -8 -3 16 105
use FILL  FILL_2090
timestamp 1711653199
transform 1 0 88 0 1 1570
box -8 -3 16 105
use FILL  FILL_2091
timestamp 1711653199
transform 1 0 80 0 1 1570
box -8 -3 16 105
use FILL  FILL_2092
timestamp 1711653199
transform 1 0 72 0 1 1570
box -8 -3 16 105
use FILL  FILL_2093
timestamp 1711653199
transform 1 0 3392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2094
timestamp 1711653199
transform 1 0 3384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2095
timestamp 1711653199
transform 1 0 3376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2096
timestamp 1711653199
transform 1 0 3344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2097
timestamp 1711653199
transform 1 0 3312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1711653199
transform 1 0 3304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1711653199
transform 1 0 3296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1711653199
transform 1 0 3288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2101
timestamp 1711653199
transform 1 0 3248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2102
timestamp 1711653199
transform 1 0 3240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2103
timestamp 1711653199
transform 1 0 3232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1711653199
transform 1 0 3192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2105
timestamp 1711653199
transform 1 0 3184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2106
timestamp 1711653199
transform 1 0 3176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1711653199
transform 1 0 3168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2108
timestamp 1711653199
transform 1 0 3160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2109
timestamp 1711653199
transform 1 0 3128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1711653199
transform 1 0 3096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1711653199
transform 1 0 3088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1711653199
transform 1 0 3048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2113
timestamp 1711653199
transform 1 0 3040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2114
timestamp 1711653199
transform 1 0 3032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2115
timestamp 1711653199
transform 1 0 2968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2116
timestamp 1711653199
transform 1 0 2960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1711653199
transform 1 0 2952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2118
timestamp 1711653199
transform 1 0 2944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2119
timestamp 1711653199
transform 1 0 2904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2120
timestamp 1711653199
transform 1 0 2896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2121
timestamp 1711653199
transform 1 0 2888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1711653199
transform 1 0 2848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2123
timestamp 1711653199
transform 1 0 2840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1711653199
transform 1 0 2832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1711653199
transform 1 0 2824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2126
timestamp 1711653199
transform 1 0 2768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2127
timestamp 1711653199
transform 1 0 2760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2128
timestamp 1711653199
transform 1 0 2752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1711653199
transform 1 0 2744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2130
timestamp 1711653199
transform 1 0 2736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2131
timestamp 1711653199
transform 1 0 2688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2132
timestamp 1711653199
transform 1 0 2680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1711653199
transform 1 0 2672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2134
timestamp 1711653199
transform 1 0 2632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1711653199
transform 1 0 2624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1711653199
transform 1 0 2616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2137
timestamp 1711653199
transform 1 0 2608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2138
timestamp 1711653199
transform 1 0 2560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2139
timestamp 1711653199
transform 1 0 2552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2140
timestamp 1711653199
transform 1 0 2544 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2141
timestamp 1711653199
transform 1 0 2536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1711653199
transform 1 0 2528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1711653199
transform 1 0 2520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2144
timestamp 1711653199
transform 1 0 2472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2145
timestamp 1711653199
transform 1 0 2464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2146
timestamp 1711653199
transform 1 0 2456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2147
timestamp 1711653199
transform 1 0 2448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2148
timestamp 1711653199
transform 1 0 2400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2149
timestamp 1711653199
transform 1 0 2392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2150
timestamp 1711653199
transform 1 0 2384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1711653199
transform 1 0 2376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1711653199
transform 1 0 2368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2153
timestamp 1711653199
transform 1 0 2360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2154
timestamp 1711653199
transform 1 0 2288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2155
timestamp 1711653199
transform 1 0 2280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1711653199
transform 1 0 2272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2157
timestamp 1711653199
transform 1 0 2264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1711653199
transform 1 0 2216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2159
timestamp 1711653199
transform 1 0 2208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1711653199
transform 1 0 2160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2161
timestamp 1711653199
transform 1 0 2152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1711653199
transform 1 0 2144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2163
timestamp 1711653199
transform 1 0 2136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2164
timestamp 1711653199
transform 1 0 2080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2165
timestamp 1711653199
transform 1 0 2072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1711653199
transform 1 0 2064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2167
timestamp 1711653199
transform 1 0 2056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1711653199
transform 1 0 1984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1711653199
transform 1 0 1976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2170
timestamp 1711653199
transform 1 0 1968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1711653199
transform 1 0 1960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2172
timestamp 1711653199
transform 1 0 1888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1711653199
transform 1 0 1880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2174
timestamp 1711653199
transform 1 0 1872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2175
timestamp 1711653199
transform 1 0 1864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2176
timestamp 1711653199
transform 1 0 1816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2177
timestamp 1711653199
transform 1 0 1792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1711653199
transform 1 0 1784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1711653199
transform 1 0 1776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2180
timestamp 1711653199
transform 1 0 1768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2181
timestamp 1711653199
transform 1 0 1744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2182
timestamp 1711653199
transform 1 0 1736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1711653199
transform 1 0 1728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2184
timestamp 1711653199
transform 1 0 1688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1711653199
transform 1 0 1680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2186
timestamp 1711653199
transform 1 0 1672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2187
timestamp 1711653199
transform 1 0 1664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1711653199
transform 1 0 1656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1711653199
transform 1 0 1608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2190
timestamp 1711653199
transform 1 0 1600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2191
timestamp 1711653199
transform 1 0 1592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1711653199
transform 1 0 1584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2193
timestamp 1711653199
transform 1 0 1576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2194
timestamp 1711653199
transform 1 0 1536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1711653199
transform 1 0 1528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2196
timestamp 1711653199
transform 1 0 1520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2197
timestamp 1711653199
transform 1 0 1512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2198
timestamp 1711653199
transform 1 0 1472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1711653199
transform 1 0 1464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2200
timestamp 1711653199
transform 1 0 1456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1711653199
transform 1 0 1448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2202
timestamp 1711653199
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1711653199
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2204
timestamp 1711653199
transform 1 0 1424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2205
timestamp 1711653199
transform 1 0 1360 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2206
timestamp 1711653199
transform 1 0 1352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2207
timestamp 1711653199
transform 1 0 1344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2208
timestamp 1711653199
transform 1 0 1336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2209
timestamp 1711653199
transform 1 0 1328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2210
timestamp 1711653199
transform 1 0 1296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2211
timestamp 1711653199
transform 1 0 1288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2212
timestamp 1711653199
transform 1 0 1280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2213
timestamp 1711653199
transform 1 0 1272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2214
timestamp 1711653199
transform 1 0 1264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2215
timestamp 1711653199
transform 1 0 1216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2216
timestamp 1711653199
transform 1 0 1208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1711653199
transform 1 0 1200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2218
timestamp 1711653199
transform 1 0 1192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2219
timestamp 1711653199
transform 1 0 1184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2220
timestamp 1711653199
transform 1 0 1176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2221
timestamp 1711653199
transform 1 0 1136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2222
timestamp 1711653199
transform 1 0 1128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2223
timestamp 1711653199
transform 1 0 1120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2224
timestamp 1711653199
transform 1 0 1112 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1711653199
transform 1 0 1072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1711653199
transform 1 0 1064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2227
timestamp 1711653199
transform 1 0 1056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2228
timestamp 1711653199
transform 1 0 1048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2229
timestamp 1711653199
transform 1 0 1040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1711653199
transform 1 0 1032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1711653199
transform 1 0 984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2232
timestamp 1711653199
transform 1 0 976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1711653199
transform 1 0 968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2234
timestamp 1711653199
transform 1 0 960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2235
timestamp 1711653199
transform 1 0 952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2236
timestamp 1711653199
transform 1 0 944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2237
timestamp 1711653199
transform 1 0 920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1711653199
transform 1 0 912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2239
timestamp 1711653199
transform 1 0 904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2240
timestamp 1711653199
transform 1 0 896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2241
timestamp 1711653199
transform 1 0 848 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2242
timestamp 1711653199
transform 1 0 840 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2243
timestamp 1711653199
transform 1 0 832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2244
timestamp 1711653199
transform 1 0 824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2245
timestamp 1711653199
transform 1 0 816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2246
timestamp 1711653199
transform 1 0 808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2247
timestamp 1711653199
transform 1 0 800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2248
timestamp 1711653199
transform 1 0 752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1711653199
transform 1 0 744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1711653199
transform 1 0 736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2251
timestamp 1711653199
transform 1 0 728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2252
timestamp 1711653199
transform 1 0 720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1711653199
transform 1 0 696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1711653199
transform 1 0 688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2255
timestamp 1711653199
transform 1 0 648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2256
timestamp 1711653199
transform 1 0 640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2257
timestamp 1711653199
transform 1 0 632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1711653199
transform 1 0 592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1711653199
transform 1 0 584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2260
timestamp 1711653199
transform 1 0 576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2261
timestamp 1711653199
transform 1 0 568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1711653199
transform 1 0 560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1711653199
transform 1 0 512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2264
timestamp 1711653199
transform 1 0 504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2265
timestamp 1711653199
transform 1 0 496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2266
timestamp 1711653199
transform 1 0 488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2267
timestamp 1711653199
transform 1 0 480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2268
timestamp 1711653199
transform 1 0 424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2269
timestamp 1711653199
transform 1 0 416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2270
timestamp 1711653199
transform 1 0 408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1711653199
transform 1 0 400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2272
timestamp 1711653199
transform 1 0 392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2273
timestamp 1711653199
transform 1 0 344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2274
timestamp 1711653199
transform 1 0 336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2275
timestamp 1711653199
transform 1 0 328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1711653199
transform 1 0 280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2277
timestamp 1711653199
transform 1 0 272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2278
timestamp 1711653199
transform 1 0 200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1711653199
transform 1 0 192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1711653199
transform 1 0 184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2281
timestamp 1711653199
transform 1 0 176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1711653199
transform 1 0 80 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2283
timestamp 1711653199
transform 1 0 72 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2284
timestamp 1711653199
transform 1 0 3392 0 1 1370
box -8 -3 16 105
use FILL  FILL_2285
timestamp 1711653199
transform 1 0 3384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2286
timestamp 1711653199
transform 1 0 3344 0 1 1370
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1711653199
transform 1 0 3336 0 1 1370
box -8 -3 16 105
use FILL  FILL_2288
timestamp 1711653199
transform 1 0 3328 0 1 1370
box -8 -3 16 105
use FILL  FILL_2289
timestamp 1711653199
transform 1 0 3320 0 1 1370
box -8 -3 16 105
use FILL  FILL_2290
timestamp 1711653199
transform 1 0 3280 0 1 1370
box -8 -3 16 105
use FILL  FILL_2291
timestamp 1711653199
transform 1 0 3272 0 1 1370
box -8 -3 16 105
use FILL  FILL_2292
timestamp 1711653199
transform 1 0 3264 0 1 1370
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1711653199
transform 1 0 3256 0 1 1370
box -8 -3 16 105
use FILL  FILL_2294
timestamp 1711653199
transform 1 0 3248 0 1 1370
box -8 -3 16 105
use FILL  FILL_2295
timestamp 1711653199
transform 1 0 3208 0 1 1370
box -8 -3 16 105
use FILL  FILL_2296
timestamp 1711653199
transform 1 0 3200 0 1 1370
box -8 -3 16 105
use FILL  FILL_2297
timestamp 1711653199
transform 1 0 3192 0 1 1370
box -8 -3 16 105
use FILL  FILL_2298
timestamp 1711653199
transform 1 0 3184 0 1 1370
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1711653199
transform 1 0 3152 0 1 1370
box -8 -3 16 105
use FILL  FILL_2300
timestamp 1711653199
transform 1 0 3144 0 1 1370
box -8 -3 16 105
use FILL  FILL_2301
timestamp 1711653199
transform 1 0 3136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1711653199
transform 1 0 3128 0 1 1370
box -8 -3 16 105
use FILL  FILL_2303
timestamp 1711653199
transform 1 0 3088 0 1 1370
box -8 -3 16 105
use FILL  FILL_2304
timestamp 1711653199
transform 1 0 3080 0 1 1370
box -8 -3 16 105
use FILL  FILL_2305
timestamp 1711653199
transform 1 0 3072 0 1 1370
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1711653199
transform 1 0 3040 0 1 1370
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1711653199
transform 1 0 3032 0 1 1370
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1711653199
transform 1 0 2992 0 1 1370
box -8 -3 16 105
use FILL  FILL_2309
timestamp 1711653199
transform 1 0 2984 0 1 1370
box -8 -3 16 105
use FILL  FILL_2310
timestamp 1711653199
transform 1 0 2976 0 1 1370
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1711653199
transform 1 0 2968 0 1 1370
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1711653199
transform 1 0 2936 0 1 1370
box -8 -3 16 105
use FILL  FILL_2313
timestamp 1711653199
transform 1 0 2928 0 1 1370
box -8 -3 16 105
use FILL  FILL_2314
timestamp 1711653199
transform 1 0 2920 0 1 1370
box -8 -3 16 105
use FILL  FILL_2315
timestamp 1711653199
transform 1 0 2888 0 1 1370
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1711653199
transform 1 0 2880 0 1 1370
box -8 -3 16 105
use FILL  FILL_2317
timestamp 1711653199
transform 1 0 2872 0 1 1370
box -8 -3 16 105
use FILL  FILL_2318
timestamp 1711653199
transform 1 0 2864 0 1 1370
box -8 -3 16 105
use FILL  FILL_2319
timestamp 1711653199
transform 1 0 2824 0 1 1370
box -8 -3 16 105
use FILL  FILL_2320
timestamp 1711653199
transform 1 0 2816 0 1 1370
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1711653199
transform 1 0 2808 0 1 1370
box -8 -3 16 105
use FILL  FILL_2322
timestamp 1711653199
transform 1 0 2800 0 1 1370
box -8 -3 16 105
use FILL  FILL_2323
timestamp 1711653199
transform 1 0 2768 0 1 1370
box -8 -3 16 105
use FILL  FILL_2324
timestamp 1711653199
transform 1 0 2760 0 1 1370
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1711653199
transform 1 0 2752 0 1 1370
box -8 -3 16 105
use FILL  FILL_2326
timestamp 1711653199
transform 1 0 2744 0 1 1370
box -8 -3 16 105
use FILL  FILL_2327
timestamp 1711653199
transform 1 0 2704 0 1 1370
box -8 -3 16 105
use FILL  FILL_2328
timestamp 1711653199
transform 1 0 2696 0 1 1370
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1711653199
transform 1 0 2656 0 1 1370
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1711653199
transform 1 0 2648 0 1 1370
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1711653199
transform 1 0 2640 0 1 1370
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1711653199
transform 1 0 2632 0 1 1370
box -8 -3 16 105
use FILL  FILL_2333
timestamp 1711653199
transform 1 0 2624 0 1 1370
box -8 -3 16 105
use FILL  FILL_2334
timestamp 1711653199
transform 1 0 2616 0 1 1370
box -8 -3 16 105
use FILL  FILL_2335
timestamp 1711653199
transform 1 0 2568 0 1 1370
box -8 -3 16 105
use FILL  FILL_2336
timestamp 1711653199
transform 1 0 2560 0 1 1370
box -8 -3 16 105
use FILL  FILL_2337
timestamp 1711653199
transform 1 0 2552 0 1 1370
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1711653199
transform 1 0 2544 0 1 1370
box -8 -3 16 105
use FILL  FILL_2339
timestamp 1711653199
transform 1 0 2536 0 1 1370
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1711653199
transform 1 0 2512 0 1 1370
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1711653199
transform 1 0 2504 0 1 1370
box -8 -3 16 105
use FILL  FILL_2342
timestamp 1711653199
transform 1 0 2472 0 1 1370
box -8 -3 16 105
use FILL  FILL_2343
timestamp 1711653199
transform 1 0 2464 0 1 1370
box -8 -3 16 105
use FILL  FILL_2344
timestamp 1711653199
transform 1 0 2456 0 1 1370
box -8 -3 16 105
use FILL  FILL_2345
timestamp 1711653199
transform 1 0 2448 0 1 1370
box -8 -3 16 105
use FILL  FILL_2346
timestamp 1711653199
transform 1 0 2416 0 1 1370
box -8 -3 16 105
use FILL  FILL_2347
timestamp 1711653199
transform 1 0 2408 0 1 1370
box -8 -3 16 105
use FILL  FILL_2348
timestamp 1711653199
transform 1 0 2384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1711653199
transform 1 0 2376 0 1 1370
box -8 -3 16 105
use FILL  FILL_2350
timestamp 1711653199
transform 1 0 2368 0 1 1370
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1711653199
transform 1 0 2328 0 1 1370
box -8 -3 16 105
use FILL  FILL_2352
timestamp 1711653199
transform 1 0 2320 0 1 1370
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1711653199
transform 1 0 2312 0 1 1370
box -8 -3 16 105
use FILL  FILL_2354
timestamp 1711653199
transform 1 0 2304 0 1 1370
box -8 -3 16 105
use FILL  FILL_2355
timestamp 1711653199
transform 1 0 2256 0 1 1370
box -8 -3 16 105
use FILL  FILL_2356
timestamp 1711653199
transform 1 0 2248 0 1 1370
box -8 -3 16 105
use FILL  FILL_2357
timestamp 1711653199
transform 1 0 2240 0 1 1370
box -8 -3 16 105
use FILL  FILL_2358
timestamp 1711653199
transform 1 0 2232 0 1 1370
box -8 -3 16 105
use FILL  FILL_2359
timestamp 1711653199
transform 1 0 2192 0 1 1370
box -8 -3 16 105
use FILL  FILL_2360
timestamp 1711653199
transform 1 0 2184 0 1 1370
box -8 -3 16 105
use FILL  FILL_2361
timestamp 1711653199
transform 1 0 2176 0 1 1370
box -8 -3 16 105
use FILL  FILL_2362
timestamp 1711653199
transform 1 0 2168 0 1 1370
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1711653199
transform 1 0 2128 0 1 1370
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1711653199
transform 1 0 2120 0 1 1370
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1711653199
transform 1 0 2112 0 1 1370
box -8 -3 16 105
use FILL  FILL_2366
timestamp 1711653199
transform 1 0 2080 0 1 1370
box -8 -3 16 105
use FILL  FILL_2367
timestamp 1711653199
transform 1 0 2072 0 1 1370
box -8 -3 16 105
use FILL  FILL_2368
timestamp 1711653199
transform 1 0 2064 0 1 1370
box -8 -3 16 105
use FILL  FILL_2369
timestamp 1711653199
transform 1 0 2056 0 1 1370
box -8 -3 16 105
use FILL  FILL_2370
timestamp 1711653199
transform 1 0 2048 0 1 1370
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1711653199
transform 1 0 1984 0 1 1370
box -8 -3 16 105
use FILL  FILL_2372
timestamp 1711653199
transform 1 0 1976 0 1 1370
box -8 -3 16 105
use FILL  FILL_2373
timestamp 1711653199
transform 1 0 1968 0 1 1370
box -8 -3 16 105
use FILL  FILL_2374
timestamp 1711653199
transform 1 0 1920 0 1 1370
box -8 -3 16 105
use FILL  FILL_2375
timestamp 1711653199
transform 1 0 1912 0 1 1370
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1711653199
transform 1 0 1904 0 1 1370
box -8 -3 16 105
use FILL  FILL_2377
timestamp 1711653199
transform 1 0 1896 0 1 1370
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1711653199
transform 1 0 1888 0 1 1370
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1711653199
transform 1 0 1848 0 1 1370
box -8 -3 16 105
use FILL  FILL_2380
timestamp 1711653199
transform 1 0 1840 0 1 1370
box -8 -3 16 105
use FILL  FILL_2381
timestamp 1711653199
transform 1 0 1832 0 1 1370
box -8 -3 16 105
use FILL  FILL_2382
timestamp 1711653199
transform 1 0 1824 0 1 1370
box -8 -3 16 105
use FILL  FILL_2383
timestamp 1711653199
transform 1 0 1816 0 1 1370
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1711653199
transform 1 0 1808 0 1 1370
box -8 -3 16 105
use FILL  FILL_2385
timestamp 1711653199
transform 1 0 1768 0 1 1370
box -8 -3 16 105
use FILL  FILL_2386
timestamp 1711653199
transform 1 0 1760 0 1 1370
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1711653199
transform 1 0 1752 0 1 1370
box -8 -3 16 105
use FILL  FILL_2388
timestamp 1711653199
transform 1 0 1744 0 1 1370
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1711653199
transform 1 0 1736 0 1 1370
box -8 -3 16 105
use FILL  FILL_2390
timestamp 1711653199
transform 1 0 1728 0 1 1370
box -8 -3 16 105
use FILL  FILL_2391
timestamp 1711653199
transform 1 0 1720 0 1 1370
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1711653199
transform 1 0 1680 0 1 1370
box -8 -3 16 105
use FILL  FILL_2393
timestamp 1711653199
transform 1 0 1672 0 1 1370
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1711653199
transform 1 0 1664 0 1 1370
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1711653199
transform 1 0 1656 0 1 1370
box -8 -3 16 105
use FILL  FILL_2396
timestamp 1711653199
transform 1 0 1624 0 1 1370
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1711653199
transform 1 0 1616 0 1 1370
box -8 -3 16 105
use FILL  FILL_2398
timestamp 1711653199
transform 1 0 1608 0 1 1370
box -8 -3 16 105
use FILL  FILL_2399
timestamp 1711653199
transform 1 0 1600 0 1 1370
box -8 -3 16 105
use FILL  FILL_2400
timestamp 1711653199
transform 1 0 1592 0 1 1370
box -8 -3 16 105
use FILL  FILL_2401
timestamp 1711653199
transform 1 0 1552 0 1 1370
box -8 -3 16 105
use FILL  FILL_2402
timestamp 1711653199
transform 1 0 1544 0 1 1370
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1711653199
transform 1 0 1536 0 1 1370
box -8 -3 16 105
use FILL  FILL_2404
timestamp 1711653199
transform 1 0 1528 0 1 1370
box -8 -3 16 105
use FILL  FILL_2405
timestamp 1711653199
transform 1 0 1520 0 1 1370
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1711653199
transform 1 0 1512 0 1 1370
box -8 -3 16 105
use FILL  FILL_2407
timestamp 1711653199
transform 1 0 1480 0 1 1370
box -8 -3 16 105
use FILL  FILL_2408
timestamp 1711653199
transform 1 0 1472 0 1 1370
box -8 -3 16 105
use FILL  FILL_2409
timestamp 1711653199
transform 1 0 1464 0 1 1370
box -8 -3 16 105
use FILL  FILL_2410
timestamp 1711653199
transform 1 0 1424 0 1 1370
box -8 -3 16 105
use FILL  FILL_2411
timestamp 1711653199
transform 1 0 1416 0 1 1370
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1711653199
transform 1 0 1408 0 1 1370
box -8 -3 16 105
use FILL  FILL_2413
timestamp 1711653199
transform 1 0 1400 0 1 1370
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1711653199
transform 1 0 1392 0 1 1370
box -8 -3 16 105
use FILL  FILL_2415
timestamp 1711653199
transform 1 0 1384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2416
timestamp 1711653199
transform 1 0 1336 0 1 1370
box -8 -3 16 105
use FILL  FILL_2417
timestamp 1711653199
transform 1 0 1328 0 1 1370
box -8 -3 16 105
use FILL  FILL_2418
timestamp 1711653199
transform 1 0 1320 0 1 1370
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1711653199
transform 1 0 1312 0 1 1370
box -8 -3 16 105
use FILL  FILL_2420
timestamp 1711653199
transform 1 0 1304 0 1 1370
box -8 -3 16 105
use FILL  FILL_2421
timestamp 1711653199
transform 1 0 1272 0 1 1370
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1711653199
transform 1 0 1240 0 1 1370
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1711653199
transform 1 0 1232 0 1 1370
box -8 -3 16 105
use FILL  FILL_2424
timestamp 1711653199
transform 1 0 1224 0 1 1370
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1711653199
transform 1 0 1216 0 1 1370
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1711653199
transform 1 0 1208 0 1 1370
box -8 -3 16 105
use FILL  FILL_2427
timestamp 1711653199
transform 1 0 1200 0 1 1370
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1711653199
transform 1 0 1192 0 1 1370
box -8 -3 16 105
use FILL  FILL_2429
timestamp 1711653199
transform 1 0 1144 0 1 1370
box -8 -3 16 105
use FILL  FILL_2430
timestamp 1711653199
transform 1 0 1136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1711653199
transform 1 0 1128 0 1 1370
box -8 -3 16 105
use FILL  FILL_2432
timestamp 1711653199
transform 1 0 1120 0 1 1370
box -8 -3 16 105
use FILL  FILL_2433
timestamp 1711653199
transform 1 0 1112 0 1 1370
box -8 -3 16 105
use FILL  FILL_2434
timestamp 1711653199
transform 1 0 1104 0 1 1370
box -8 -3 16 105
use FILL  FILL_2435
timestamp 1711653199
transform 1 0 1064 0 1 1370
box -8 -3 16 105
use FILL  FILL_2436
timestamp 1711653199
transform 1 0 1056 0 1 1370
box -8 -3 16 105
use FILL  FILL_2437
timestamp 1711653199
transform 1 0 1048 0 1 1370
box -8 -3 16 105
use FILL  FILL_2438
timestamp 1711653199
transform 1 0 1040 0 1 1370
box -8 -3 16 105
use FILL  FILL_2439
timestamp 1711653199
transform 1 0 1008 0 1 1370
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1711653199
transform 1 0 1000 0 1 1370
box -8 -3 16 105
use FILL  FILL_2441
timestamp 1711653199
transform 1 0 992 0 1 1370
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1711653199
transform 1 0 984 0 1 1370
box -8 -3 16 105
use FILL  FILL_2443
timestamp 1711653199
transform 1 0 976 0 1 1370
box -8 -3 16 105
use FILL  FILL_2444
timestamp 1711653199
transform 1 0 936 0 1 1370
box -8 -3 16 105
use FILL  FILL_2445
timestamp 1711653199
transform 1 0 928 0 1 1370
box -8 -3 16 105
use FILL  FILL_2446
timestamp 1711653199
transform 1 0 920 0 1 1370
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1711653199
transform 1 0 880 0 1 1370
box -8 -3 16 105
use FILL  FILL_2448
timestamp 1711653199
transform 1 0 872 0 1 1370
box -8 -3 16 105
use FILL  FILL_2449
timestamp 1711653199
transform 1 0 864 0 1 1370
box -8 -3 16 105
use FILL  FILL_2450
timestamp 1711653199
transform 1 0 856 0 1 1370
box -8 -3 16 105
use FILL  FILL_2451
timestamp 1711653199
transform 1 0 848 0 1 1370
box -8 -3 16 105
use FILL  FILL_2452
timestamp 1711653199
transform 1 0 816 0 1 1370
box -8 -3 16 105
use FILL  FILL_2453
timestamp 1711653199
transform 1 0 808 0 1 1370
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1711653199
transform 1 0 800 0 1 1370
box -8 -3 16 105
use FILL  FILL_2455
timestamp 1711653199
transform 1 0 792 0 1 1370
box -8 -3 16 105
use FILL  FILL_2456
timestamp 1711653199
transform 1 0 744 0 1 1370
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1711653199
transform 1 0 736 0 1 1370
box -8 -3 16 105
use FILL  FILL_2458
timestamp 1711653199
transform 1 0 728 0 1 1370
box -8 -3 16 105
use FILL  FILL_2459
timestamp 1711653199
transform 1 0 720 0 1 1370
box -8 -3 16 105
use FILL  FILL_2460
timestamp 1711653199
transform 1 0 672 0 1 1370
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1711653199
transform 1 0 664 0 1 1370
box -8 -3 16 105
use FILL  FILL_2462
timestamp 1711653199
transform 1 0 656 0 1 1370
box -8 -3 16 105
use FILL  FILL_2463
timestamp 1711653199
transform 1 0 608 0 1 1370
box -8 -3 16 105
use FILL  FILL_2464
timestamp 1711653199
transform 1 0 600 0 1 1370
box -8 -3 16 105
use FILL  FILL_2465
timestamp 1711653199
transform 1 0 592 0 1 1370
box -8 -3 16 105
use FILL  FILL_2466
timestamp 1711653199
transform 1 0 584 0 1 1370
box -8 -3 16 105
use FILL  FILL_2467
timestamp 1711653199
transform 1 0 544 0 1 1370
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1711653199
transform 1 0 536 0 1 1370
box -8 -3 16 105
use FILL  FILL_2469
timestamp 1711653199
transform 1 0 488 0 1 1370
box -8 -3 16 105
use FILL  FILL_2470
timestamp 1711653199
transform 1 0 480 0 1 1370
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1711653199
transform 1 0 472 0 1 1370
box -8 -3 16 105
use FILL  FILL_2472
timestamp 1711653199
transform 1 0 464 0 1 1370
box -8 -3 16 105
use FILL  FILL_2473
timestamp 1711653199
transform 1 0 392 0 1 1370
box -8 -3 16 105
use FILL  FILL_2474
timestamp 1711653199
transform 1 0 384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1711653199
transform 1 0 376 0 1 1370
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1711653199
transform 1 0 328 0 1 1370
box -8 -3 16 105
use FILL  FILL_2477
timestamp 1711653199
transform 1 0 280 0 1 1370
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1711653199
transform 1 0 272 0 1 1370
box -8 -3 16 105
use FILL  FILL_2479
timestamp 1711653199
transform 1 0 264 0 1 1370
box -8 -3 16 105
use FILL  FILL_2480
timestamp 1711653199
transform 1 0 256 0 1 1370
box -8 -3 16 105
use FILL  FILL_2481
timestamp 1711653199
transform 1 0 248 0 1 1370
box -8 -3 16 105
use FILL  FILL_2482
timestamp 1711653199
transform 1 0 184 0 1 1370
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1711653199
transform 1 0 176 0 1 1370
box -8 -3 16 105
use FILL  FILL_2484
timestamp 1711653199
transform 1 0 168 0 1 1370
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1711653199
transform 1 0 128 0 1 1370
box -8 -3 16 105
use FILL  FILL_2486
timestamp 1711653199
transform 1 0 120 0 1 1370
box -8 -3 16 105
use FILL  FILL_2487
timestamp 1711653199
transform 1 0 80 0 1 1370
box -8 -3 16 105
use FILL  FILL_2488
timestamp 1711653199
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_2489
timestamp 1711653199
transform 1 0 3392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2490
timestamp 1711653199
transform 1 0 3384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2491
timestamp 1711653199
transform 1 0 3344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1711653199
transform 1 0 3336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2493
timestamp 1711653199
transform 1 0 3328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1711653199
transform 1 0 3288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2495
timestamp 1711653199
transform 1 0 3280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2496
timestamp 1711653199
transform 1 0 3272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2497
timestamp 1711653199
transform 1 0 3264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2498
timestamp 1711653199
transform 1 0 3232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2499
timestamp 1711653199
transform 1 0 3224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1711653199
transform 1 0 3192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1711653199
transform 1 0 3184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2502
timestamp 1711653199
transform 1 0 3176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2503
timestamp 1711653199
transform 1 0 3168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2504
timestamp 1711653199
transform 1 0 3128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2505
timestamp 1711653199
transform 1 0 3120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1711653199
transform 1 0 3112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2507
timestamp 1711653199
transform 1 0 3072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1711653199
transform 1 0 3064 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2509
timestamp 1711653199
transform 1 0 3056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1711653199
transform 1 0 3048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1711653199
transform 1 0 3040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2512
timestamp 1711653199
transform 1 0 3032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2513
timestamp 1711653199
transform 1 0 2976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1711653199
transform 1 0 2968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2515
timestamp 1711653199
transform 1 0 2960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2516
timestamp 1711653199
transform 1 0 2952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2517
timestamp 1711653199
transform 1 0 2944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2518
timestamp 1711653199
transform 1 0 2904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1711653199
transform 1 0 2896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2520
timestamp 1711653199
transform 1 0 2856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2521
timestamp 1711653199
transform 1 0 2848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1711653199
transform 1 0 2840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1711653199
transform 1 0 2832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2524
timestamp 1711653199
transform 1 0 2792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1711653199
transform 1 0 2784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2526
timestamp 1711653199
transform 1 0 2776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1711653199
transform 1 0 2768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2528
timestamp 1711653199
transform 1 0 2728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1711653199
transform 1 0 2720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1711653199
transform 1 0 2680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2531
timestamp 1711653199
transform 1 0 2672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2532
timestamp 1711653199
transform 1 0 2664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2533
timestamp 1711653199
transform 1 0 2632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1711653199
transform 1 0 2624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2535
timestamp 1711653199
transform 1 0 2616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2536
timestamp 1711653199
transform 1 0 2608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2537
timestamp 1711653199
transform 1 0 2560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1711653199
transform 1 0 2552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1711653199
transform 1 0 2544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2540
timestamp 1711653199
transform 1 0 2536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1711653199
transform 1 0 2488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2542
timestamp 1711653199
transform 1 0 2480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1711653199
transform 1 0 2472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2544
timestamp 1711653199
transform 1 0 2464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1711653199
transform 1 0 2456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2546
timestamp 1711653199
transform 1 0 2408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1711653199
transform 1 0 2400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2548
timestamp 1711653199
transform 1 0 2392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2549
timestamp 1711653199
transform 1 0 2360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2550
timestamp 1711653199
transform 1 0 2352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2551
timestamp 1711653199
transform 1 0 2344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2552
timestamp 1711653199
transform 1 0 2320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2553
timestamp 1711653199
transform 1 0 2312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1711653199
transform 1 0 2304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2555
timestamp 1711653199
transform 1 0 2272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1711653199
transform 1 0 2264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2557
timestamp 1711653199
transform 1 0 2256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1711653199
transform 1 0 2248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2559
timestamp 1711653199
transform 1 0 2208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2560
timestamp 1711653199
transform 1 0 2200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1711653199
transform 1 0 2192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2562
timestamp 1711653199
transform 1 0 2184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2563
timestamp 1711653199
transform 1 0 2136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2564
timestamp 1711653199
transform 1 0 2128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2565
timestamp 1711653199
transform 1 0 2120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2566
timestamp 1711653199
transform 1 0 2112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2567
timestamp 1711653199
transform 1 0 2104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1711653199
transform 1 0 2096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1711653199
transform 1 0 2048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2570
timestamp 1711653199
transform 1 0 2040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2571
timestamp 1711653199
transform 1 0 2032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2572
timestamp 1711653199
transform 1 0 1992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1711653199
transform 1 0 1984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2574
timestamp 1711653199
transform 1 0 1976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2575
timestamp 1711653199
transform 1 0 1968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2576
timestamp 1711653199
transform 1 0 1936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2577
timestamp 1711653199
transform 1 0 1928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2578
timestamp 1711653199
transform 1 0 1920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2579
timestamp 1711653199
transform 1 0 1872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1711653199
transform 1 0 1864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2581
timestamp 1711653199
transform 1 0 1856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2582
timestamp 1711653199
transform 1 0 1848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2583
timestamp 1711653199
transform 1 0 1840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1711653199
transform 1 0 1808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1711653199
transform 1 0 1800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2586
timestamp 1711653199
transform 1 0 1792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2587
timestamp 1711653199
transform 1 0 1784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2588
timestamp 1711653199
transform 1 0 1776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2589
timestamp 1711653199
transform 1 0 1728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2590
timestamp 1711653199
transform 1 0 1720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1711653199
transform 1 0 1712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2592
timestamp 1711653199
transform 1 0 1704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1711653199
transform 1 0 1696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1711653199
transform 1 0 1688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2595
timestamp 1711653199
transform 1 0 1680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2596
timestamp 1711653199
transform 1 0 1648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1711653199
transform 1 0 1640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1711653199
transform 1 0 1632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2599
timestamp 1711653199
transform 1 0 1624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2600
timestamp 1711653199
transform 1 0 1584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2601
timestamp 1711653199
transform 1 0 1576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2602
timestamp 1711653199
transform 1 0 1568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2603
timestamp 1711653199
transform 1 0 1560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2604
timestamp 1711653199
transform 1 0 1552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1711653199
transform 1 0 1544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2606
timestamp 1711653199
transform 1 0 1536 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2607
timestamp 1711653199
transform 1 0 1496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1711653199
transform 1 0 1488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2609
timestamp 1711653199
transform 1 0 1480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2610
timestamp 1711653199
transform 1 0 1472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2611
timestamp 1711653199
transform 1 0 1464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2612
timestamp 1711653199
transform 1 0 1456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2613
timestamp 1711653199
transform 1 0 1424 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1711653199
transform 1 0 1416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2615
timestamp 1711653199
transform 1 0 1408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2616
timestamp 1711653199
transform 1 0 1400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2617
timestamp 1711653199
transform 1 0 1368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2618
timestamp 1711653199
transform 1 0 1360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2619
timestamp 1711653199
transform 1 0 1352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1711653199
transform 1 0 1344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2621
timestamp 1711653199
transform 1 0 1336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2622
timestamp 1711653199
transform 1 0 1328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1711653199
transform 1 0 1288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2624
timestamp 1711653199
transform 1 0 1280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2625
timestamp 1711653199
transform 1 0 1272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1711653199
transform 1 0 1264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2627
timestamp 1711653199
transform 1 0 1256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2628
timestamp 1711653199
transform 1 0 1248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1711653199
transform 1 0 1208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2630
timestamp 1711653199
transform 1 0 1200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2631
timestamp 1711653199
transform 1 0 1192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2632
timestamp 1711653199
transform 1 0 1184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1711653199
transform 1 0 1176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2634
timestamp 1711653199
transform 1 0 1168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2635
timestamp 1711653199
transform 1 0 1128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2636
timestamp 1711653199
transform 1 0 1120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2637
timestamp 1711653199
transform 1 0 1112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2638
timestamp 1711653199
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2639
timestamp 1711653199
transform 1 0 1096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2640
timestamp 1711653199
transform 1 0 1056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2641
timestamp 1711653199
transform 1 0 1048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2642
timestamp 1711653199
transform 1 0 1040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2643
timestamp 1711653199
transform 1 0 1032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1711653199
transform 1 0 992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1711653199
transform 1 0 984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2646
timestamp 1711653199
transform 1 0 976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2647
timestamp 1711653199
transform 1 0 968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1711653199
transform 1 0 960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2649
timestamp 1711653199
transform 1 0 920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1711653199
transform 1 0 912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2651
timestamp 1711653199
transform 1 0 904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2652
timestamp 1711653199
transform 1 0 896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1711653199
transform 1 0 856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2654
timestamp 1711653199
transform 1 0 848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1711653199
transform 1 0 840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2656
timestamp 1711653199
transform 1 0 800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2657
timestamp 1711653199
transform 1 0 792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1711653199
transform 1 0 784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2659
timestamp 1711653199
transform 1 0 776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2660
timestamp 1711653199
transform 1 0 736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1711653199
transform 1 0 712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2662
timestamp 1711653199
transform 1 0 704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2663
timestamp 1711653199
transform 1 0 696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2664
timestamp 1711653199
transform 1 0 688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1711653199
transform 1 0 648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1711653199
transform 1 0 640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2667
timestamp 1711653199
transform 1 0 592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1711653199
transform 1 0 584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2669
timestamp 1711653199
transform 1 0 576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1711653199
transform 1 0 568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2671
timestamp 1711653199
transform 1 0 560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2672
timestamp 1711653199
transform 1 0 552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1711653199
transform 1 0 544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2674
timestamp 1711653199
transform 1 0 480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2675
timestamp 1711653199
transform 1 0 472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2676
timestamp 1711653199
transform 1 0 464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2677
timestamp 1711653199
transform 1 0 456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2678
timestamp 1711653199
transform 1 0 448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1711653199
transform 1 0 440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1711653199
transform 1 0 376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2681
timestamp 1711653199
transform 1 0 368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2682
timestamp 1711653199
transform 1 0 360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1711653199
transform 1 0 352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2684
timestamp 1711653199
transform 1 0 344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2685
timestamp 1711653199
transform 1 0 336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2686
timestamp 1711653199
transform 1 0 328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2687
timestamp 1711653199
transform 1 0 280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2688
timestamp 1711653199
transform 1 0 272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2689
timestamp 1711653199
transform 1 0 264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1711653199
transform 1 0 224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2691
timestamp 1711653199
transform 1 0 216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2692
timestamp 1711653199
transform 1 0 208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1711653199
transform 1 0 200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2694
timestamp 1711653199
transform 1 0 192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2695
timestamp 1711653199
transform 1 0 184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2696
timestamp 1711653199
transform 1 0 136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2697
timestamp 1711653199
transform 1 0 128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1711653199
transform 1 0 120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1711653199
transform 1 0 112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2700
timestamp 1711653199
transform 1 0 80 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2701
timestamp 1711653199
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2702
timestamp 1711653199
transform 1 0 3392 0 1 1170
box -8 -3 16 105
use FILL  FILL_2703
timestamp 1711653199
transform 1 0 3384 0 1 1170
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1711653199
transform 1 0 3376 0 1 1170
box -8 -3 16 105
use FILL  FILL_2705
timestamp 1711653199
transform 1 0 3328 0 1 1170
box -8 -3 16 105
use FILL  FILL_2706
timestamp 1711653199
transform 1 0 3320 0 1 1170
box -8 -3 16 105
use FILL  FILL_2707
timestamp 1711653199
transform 1 0 3312 0 1 1170
box -8 -3 16 105
use FILL  FILL_2708
timestamp 1711653199
transform 1 0 3304 0 1 1170
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1711653199
transform 1 0 3296 0 1 1170
box -8 -3 16 105
use FILL  FILL_2710
timestamp 1711653199
transform 1 0 3248 0 1 1170
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1711653199
transform 1 0 3240 0 1 1170
box -8 -3 16 105
use FILL  FILL_2712
timestamp 1711653199
transform 1 0 3232 0 1 1170
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1711653199
transform 1 0 3224 0 1 1170
box -8 -3 16 105
use FILL  FILL_2714
timestamp 1711653199
transform 1 0 3216 0 1 1170
box -8 -3 16 105
use FILL  FILL_2715
timestamp 1711653199
transform 1 0 3176 0 1 1170
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1711653199
transform 1 0 3168 0 1 1170
box -8 -3 16 105
use FILL  FILL_2717
timestamp 1711653199
transform 1 0 3160 0 1 1170
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1711653199
transform 1 0 3152 0 1 1170
box -8 -3 16 105
use FILL  FILL_2719
timestamp 1711653199
transform 1 0 3144 0 1 1170
box -8 -3 16 105
use FILL  FILL_2720
timestamp 1711653199
transform 1 0 3096 0 1 1170
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1711653199
transform 1 0 3088 0 1 1170
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1711653199
transform 1 0 3080 0 1 1170
box -8 -3 16 105
use FILL  FILL_2723
timestamp 1711653199
transform 1 0 3072 0 1 1170
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1711653199
transform 1 0 3064 0 1 1170
box -8 -3 16 105
use FILL  FILL_2725
timestamp 1711653199
transform 1 0 3024 0 1 1170
box -8 -3 16 105
use FILL  FILL_2726
timestamp 1711653199
transform 1 0 3016 0 1 1170
box -8 -3 16 105
use FILL  FILL_2727
timestamp 1711653199
transform 1 0 2976 0 1 1170
box -8 -3 16 105
use FILL  FILL_2728
timestamp 1711653199
transform 1 0 2968 0 1 1170
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1711653199
transform 1 0 2960 0 1 1170
box -8 -3 16 105
use FILL  FILL_2730
timestamp 1711653199
transform 1 0 2952 0 1 1170
box -8 -3 16 105
use FILL  FILL_2731
timestamp 1711653199
transform 1 0 2944 0 1 1170
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1711653199
transform 1 0 2936 0 1 1170
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1711653199
transform 1 0 2880 0 1 1170
box -8 -3 16 105
use FILL  FILL_2734
timestamp 1711653199
transform 1 0 2872 0 1 1170
box -8 -3 16 105
use FILL  FILL_2735
timestamp 1711653199
transform 1 0 2864 0 1 1170
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1711653199
transform 1 0 2856 0 1 1170
box -8 -3 16 105
use FILL  FILL_2737
timestamp 1711653199
transform 1 0 2848 0 1 1170
box -8 -3 16 105
use FILL  FILL_2738
timestamp 1711653199
transform 1 0 2800 0 1 1170
box -8 -3 16 105
use FILL  FILL_2739
timestamp 1711653199
transform 1 0 2792 0 1 1170
box -8 -3 16 105
use FILL  FILL_2740
timestamp 1711653199
transform 1 0 2784 0 1 1170
box -8 -3 16 105
use FILL  FILL_2741
timestamp 1711653199
transform 1 0 2776 0 1 1170
box -8 -3 16 105
use FILL  FILL_2742
timestamp 1711653199
transform 1 0 2736 0 1 1170
box -8 -3 16 105
use FILL  FILL_2743
timestamp 1711653199
transform 1 0 2728 0 1 1170
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1711653199
transform 1 0 2720 0 1 1170
box -8 -3 16 105
use FILL  FILL_2745
timestamp 1711653199
transform 1 0 2672 0 1 1170
box -8 -3 16 105
use FILL  FILL_2746
timestamp 1711653199
transform 1 0 2664 0 1 1170
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1711653199
transform 1 0 2656 0 1 1170
box -8 -3 16 105
use FILL  FILL_2748
timestamp 1711653199
transform 1 0 2648 0 1 1170
box -8 -3 16 105
use FILL  FILL_2749
timestamp 1711653199
transform 1 0 2640 0 1 1170
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1711653199
transform 1 0 2592 0 1 1170
box -8 -3 16 105
use FILL  FILL_2751
timestamp 1711653199
transform 1 0 2584 0 1 1170
box -8 -3 16 105
use FILL  FILL_2752
timestamp 1711653199
transform 1 0 2576 0 1 1170
box -8 -3 16 105
use FILL  FILL_2753
timestamp 1711653199
transform 1 0 2552 0 1 1170
box -8 -3 16 105
use FILL  FILL_2754
timestamp 1711653199
transform 1 0 2544 0 1 1170
box -8 -3 16 105
use FILL  FILL_2755
timestamp 1711653199
transform 1 0 2536 0 1 1170
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1711653199
transform 1 0 2504 0 1 1170
box -8 -3 16 105
use FILL  FILL_2757
timestamp 1711653199
transform 1 0 2496 0 1 1170
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1711653199
transform 1 0 2456 0 1 1170
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1711653199
transform 1 0 2448 0 1 1170
box -8 -3 16 105
use FILL  FILL_2760
timestamp 1711653199
transform 1 0 2440 0 1 1170
box -8 -3 16 105
use FILL  FILL_2761
timestamp 1711653199
transform 1 0 2432 0 1 1170
box -8 -3 16 105
use FILL  FILL_2762
timestamp 1711653199
transform 1 0 2424 0 1 1170
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1711653199
transform 1 0 2368 0 1 1170
box -8 -3 16 105
use FILL  FILL_2764
timestamp 1711653199
transform 1 0 2360 0 1 1170
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1711653199
transform 1 0 2352 0 1 1170
box -8 -3 16 105
use FILL  FILL_2766
timestamp 1711653199
transform 1 0 2328 0 1 1170
box -8 -3 16 105
use FILL  FILL_2767
timestamp 1711653199
transform 1 0 2320 0 1 1170
box -8 -3 16 105
use FILL  FILL_2768
timestamp 1711653199
transform 1 0 2312 0 1 1170
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1711653199
transform 1 0 2304 0 1 1170
box -8 -3 16 105
use FILL  FILL_2770
timestamp 1711653199
transform 1 0 2264 0 1 1170
box -8 -3 16 105
use FILL  FILL_2771
timestamp 1711653199
transform 1 0 2256 0 1 1170
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1711653199
transform 1 0 2248 0 1 1170
box -8 -3 16 105
use FILL  FILL_2773
timestamp 1711653199
transform 1 0 2240 0 1 1170
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1711653199
transform 1 0 2200 0 1 1170
box -8 -3 16 105
use FILL  FILL_2775
timestamp 1711653199
transform 1 0 2192 0 1 1170
box -8 -3 16 105
use FILL  FILL_2776
timestamp 1711653199
transform 1 0 2184 0 1 1170
box -8 -3 16 105
use FILL  FILL_2777
timestamp 1711653199
transform 1 0 2176 0 1 1170
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1711653199
transform 1 0 2168 0 1 1170
box -8 -3 16 105
use FILL  FILL_2779
timestamp 1711653199
transform 1 0 2128 0 1 1170
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1711653199
transform 1 0 2120 0 1 1170
box -8 -3 16 105
use FILL  FILL_2781
timestamp 1711653199
transform 1 0 2112 0 1 1170
box -8 -3 16 105
use FILL  FILL_2782
timestamp 1711653199
transform 1 0 2104 0 1 1170
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1711653199
transform 1 0 2096 0 1 1170
box -8 -3 16 105
use FILL  FILL_2784
timestamp 1711653199
transform 1 0 2072 0 1 1170
box -8 -3 16 105
use FILL  FILL_2785
timestamp 1711653199
transform 1 0 2040 0 1 1170
box -8 -3 16 105
use FILL  FILL_2786
timestamp 1711653199
transform 1 0 2032 0 1 1170
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1711653199
transform 1 0 2024 0 1 1170
box -8 -3 16 105
use FILL  FILL_2788
timestamp 1711653199
transform 1 0 2016 0 1 1170
box -8 -3 16 105
use FILL  FILL_2789
timestamp 1711653199
transform 1 0 2008 0 1 1170
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1711653199
transform 1 0 2000 0 1 1170
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1711653199
transform 1 0 1952 0 1 1170
box -8 -3 16 105
use FILL  FILL_2792
timestamp 1711653199
transform 1 0 1944 0 1 1170
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1711653199
transform 1 0 1936 0 1 1170
box -8 -3 16 105
use FILL  FILL_2794
timestamp 1711653199
transform 1 0 1928 0 1 1170
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1711653199
transform 1 0 1888 0 1 1170
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1711653199
transform 1 0 1880 0 1 1170
box -8 -3 16 105
use FILL  FILL_2797
timestamp 1711653199
transform 1 0 1872 0 1 1170
box -8 -3 16 105
use FILL  FILL_2798
timestamp 1711653199
transform 1 0 1864 0 1 1170
box -8 -3 16 105
use FILL  FILL_2799
timestamp 1711653199
transform 1 0 1856 0 1 1170
box -8 -3 16 105
use FILL  FILL_2800
timestamp 1711653199
transform 1 0 1848 0 1 1170
box -8 -3 16 105
use FILL  FILL_2801
timestamp 1711653199
transform 1 0 1808 0 1 1170
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1711653199
transform 1 0 1800 0 1 1170
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1711653199
transform 1 0 1792 0 1 1170
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1711653199
transform 1 0 1784 0 1 1170
box -8 -3 16 105
use FILL  FILL_2805
timestamp 1711653199
transform 1 0 1776 0 1 1170
box -8 -3 16 105
use FILL  FILL_2806
timestamp 1711653199
transform 1 0 1768 0 1 1170
box -8 -3 16 105
use FILL  FILL_2807
timestamp 1711653199
transform 1 0 1728 0 1 1170
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1711653199
transform 1 0 1720 0 1 1170
box -8 -3 16 105
use FILL  FILL_2809
timestamp 1711653199
transform 1 0 1712 0 1 1170
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1711653199
transform 1 0 1704 0 1 1170
box -8 -3 16 105
use FILL  FILL_2811
timestamp 1711653199
transform 1 0 1696 0 1 1170
box -8 -3 16 105
use FILL  FILL_2812
timestamp 1711653199
transform 1 0 1688 0 1 1170
box -8 -3 16 105
use FILL  FILL_2813
timestamp 1711653199
transform 1 0 1680 0 1 1170
box -8 -3 16 105
use FILL  FILL_2814
timestamp 1711653199
transform 1 0 1672 0 1 1170
box -8 -3 16 105
use FILL  FILL_2815
timestamp 1711653199
transform 1 0 1624 0 1 1170
box -8 -3 16 105
use FILL  FILL_2816
timestamp 1711653199
transform 1 0 1616 0 1 1170
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1711653199
transform 1 0 1608 0 1 1170
box -8 -3 16 105
use FILL  FILL_2818
timestamp 1711653199
transform 1 0 1600 0 1 1170
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1711653199
transform 1 0 1592 0 1 1170
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1711653199
transform 1 0 1584 0 1 1170
box -8 -3 16 105
use FILL  FILL_2821
timestamp 1711653199
transform 1 0 1576 0 1 1170
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1711653199
transform 1 0 1568 0 1 1170
box -8 -3 16 105
use FILL  FILL_2823
timestamp 1711653199
transform 1 0 1528 0 1 1170
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1711653199
transform 1 0 1520 0 1 1170
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1711653199
transform 1 0 1512 0 1 1170
box -8 -3 16 105
use FILL  FILL_2826
timestamp 1711653199
transform 1 0 1504 0 1 1170
box -8 -3 16 105
use FILL  FILL_2827
timestamp 1711653199
transform 1 0 1496 0 1 1170
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1711653199
transform 1 0 1456 0 1 1170
box -8 -3 16 105
use FILL  FILL_2829
timestamp 1711653199
transform 1 0 1448 0 1 1170
box -8 -3 16 105
use FILL  FILL_2830
timestamp 1711653199
transform 1 0 1440 0 1 1170
box -8 -3 16 105
use FILL  FILL_2831
timestamp 1711653199
transform 1 0 1432 0 1 1170
box -8 -3 16 105
use FILL  FILL_2832
timestamp 1711653199
transform 1 0 1424 0 1 1170
box -8 -3 16 105
use FILL  FILL_2833
timestamp 1711653199
transform 1 0 1392 0 1 1170
box -8 -3 16 105
use FILL  FILL_2834
timestamp 1711653199
transform 1 0 1384 0 1 1170
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1711653199
transform 1 0 1376 0 1 1170
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1711653199
transform 1 0 1368 0 1 1170
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1711653199
transform 1 0 1360 0 1 1170
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1711653199
transform 1 0 1352 0 1 1170
box -8 -3 16 105
use FILL  FILL_2839
timestamp 1711653199
transform 1 0 1312 0 1 1170
box -8 -3 16 105
use FILL  FILL_2840
timestamp 1711653199
transform 1 0 1304 0 1 1170
box -8 -3 16 105
use FILL  FILL_2841
timestamp 1711653199
transform 1 0 1296 0 1 1170
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1711653199
transform 1 0 1288 0 1 1170
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1711653199
transform 1 0 1280 0 1 1170
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1711653199
transform 1 0 1272 0 1 1170
box -8 -3 16 105
use FILL  FILL_2845
timestamp 1711653199
transform 1 0 1264 0 1 1170
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1711653199
transform 1 0 1256 0 1 1170
box -8 -3 16 105
use FILL  FILL_2847
timestamp 1711653199
transform 1 0 1248 0 1 1170
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1711653199
transform 1 0 1200 0 1 1170
box -8 -3 16 105
use FILL  FILL_2849
timestamp 1711653199
transform 1 0 1192 0 1 1170
box -8 -3 16 105
use FILL  FILL_2850
timestamp 1711653199
transform 1 0 1184 0 1 1170
box -8 -3 16 105
use FILL  FILL_2851
timestamp 1711653199
transform 1 0 1176 0 1 1170
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1711653199
transform 1 0 1168 0 1 1170
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1711653199
transform 1 0 1160 0 1 1170
box -8 -3 16 105
use FILL  FILL_2854
timestamp 1711653199
transform 1 0 1152 0 1 1170
box -8 -3 16 105
use FILL  FILL_2855
timestamp 1711653199
transform 1 0 1144 0 1 1170
box -8 -3 16 105
use FILL  FILL_2856
timestamp 1711653199
transform 1 0 1120 0 1 1170
box -8 -3 16 105
use FILL  FILL_2857
timestamp 1711653199
transform 1 0 1112 0 1 1170
box -8 -3 16 105
use FILL  FILL_2858
timestamp 1711653199
transform 1 0 1072 0 1 1170
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1711653199
transform 1 0 1064 0 1 1170
box -8 -3 16 105
use FILL  FILL_2860
timestamp 1711653199
transform 1 0 1056 0 1 1170
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1711653199
transform 1 0 1048 0 1 1170
box -8 -3 16 105
use FILL  FILL_2862
timestamp 1711653199
transform 1 0 1040 0 1 1170
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1711653199
transform 1 0 1032 0 1 1170
box -8 -3 16 105
use FILL  FILL_2864
timestamp 1711653199
transform 1 0 1024 0 1 1170
box -8 -3 16 105
use FILL  FILL_2865
timestamp 1711653199
transform 1 0 1016 0 1 1170
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1711653199
transform 1 0 968 0 1 1170
box -8 -3 16 105
use FILL  FILL_2867
timestamp 1711653199
transform 1 0 960 0 1 1170
box -8 -3 16 105
use FILL  FILL_2868
timestamp 1711653199
transform 1 0 952 0 1 1170
box -8 -3 16 105
use FILL  FILL_2869
timestamp 1711653199
transform 1 0 944 0 1 1170
box -8 -3 16 105
use FILL  FILL_2870
timestamp 1711653199
transform 1 0 936 0 1 1170
box -8 -3 16 105
use FILL  FILL_2871
timestamp 1711653199
transform 1 0 928 0 1 1170
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1711653199
transform 1 0 920 0 1 1170
box -8 -3 16 105
use FILL  FILL_2873
timestamp 1711653199
transform 1 0 912 0 1 1170
box -8 -3 16 105
use FILL  FILL_2874
timestamp 1711653199
transform 1 0 872 0 1 1170
box -8 -3 16 105
use FILL  FILL_2875
timestamp 1711653199
transform 1 0 864 0 1 1170
box -8 -3 16 105
use FILL  FILL_2876
timestamp 1711653199
transform 1 0 856 0 1 1170
box -8 -3 16 105
use FILL  FILL_2877
timestamp 1711653199
transform 1 0 848 0 1 1170
box -8 -3 16 105
use FILL  FILL_2878
timestamp 1711653199
transform 1 0 840 0 1 1170
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1711653199
transform 1 0 832 0 1 1170
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1711653199
transform 1 0 792 0 1 1170
box -8 -3 16 105
use FILL  FILL_2881
timestamp 1711653199
transform 1 0 784 0 1 1170
box -8 -3 16 105
use FILL  FILL_2882
timestamp 1711653199
transform 1 0 776 0 1 1170
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1711653199
transform 1 0 768 0 1 1170
box -8 -3 16 105
use FILL  FILL_2884
timestamp 1711653199
transform 1 0 728 0 1 1170
box -8 -3 16 105
use FILL  FILL_2885
timestamp 1711653199
transform 1 0 720 0 1 1170
box -8 -3 16 105
use FILL  FILL_2886
timestamp 1711653199
transform 1 0 712 0 1 1170
box -8 -3 16 105
use FILL  FILL_2887
timestamp 1711653199
transform 1 0 704 0 1 1170
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1711653199
transform 1 0 672 0 1 1170
box -8 -3 16 105
use FILL  FILL_2889
timestamp 1711653199
transform 1 0 664 0 1 1170
box -8 -3 16 105
use FILL  FILL_2890
timestamp 1711653199
transform 1 0 656 0 1 1170
box -8 -3 16 105
use FILL  FILL_2891
timestamp 1711653199
transform 1 0 648 0 1 1170
box -8 -3 16 105
use FILL  FILL_2892
timestamp 1711653199
transform 1 0 616 0 1 1170
box -8 -3 16 105
use FILL  FILL_2893
timestamp 1711653199
transform 1 0 608 0 1 1170
box -8 -3 16 105
use FILL  FILL_2894
timestamp 1711653199
transform 1 0 600 0 1 1170
box -8 -3 16 105
use FILL  FILL_2895
timestamp 1711653199
transform 1 0 568 0 1 1170
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1711653199
transform 1 0 560 0 1 1170
box -8 -3 16 105
use FILL  FILL_2897
timestamp 1711653199
transform 1 0 552 0 1 1170
box -8 -3 16 105
use FILL  FILL_2898
timestamp 1711653199
transform 1 0 544 0 1 1170
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1711653199
transform 1 0 504 0 1 1170
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1711653199
transform 1 0 496 0 1 1170
box -8 -3 16 105
use FILL  FILL_2901
timestamp 1711653199
transform 1 0 488 0 1 1170
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1711653199
transform 1 0 480 0 1 1170
box -8 -3 16 105
use FILL  FILL_2903
timestamp 1711653199
transform 1 0 440 0 1 1170
box -8 -3 16 105
use FILL  FILL_2904
timestamp 1711653199
transform 1 0 432 0 1 1170
box -8 -3 16 105
use FILL  FILL_2905
timestamp 1711653199
transform 1 0 424 0 1 1170
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1711653199
transform 1 0 392 0 1 1170
box -8 -3 16 105
use FILL  FILL_2907
timestamp 1711653199
transform 1 0 384 0 1 1170
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1711653199
transform 1 0 376 0 1 1170
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1711653199
transform 1 0 344 0 1 1170
box -8 -3 16 105
use FILL  FILL_2910
timestamp 1711653199
transform 1 0 336 0 1 1170
box -8 -3 16 105
use FILL  FILL_2911
timestamp 1711653199
transform 1 0 328 0 1 1170
box -8 -3 16 105
use FILL  FILL_2912
timestamp 1711653199
transform 1 0 320 0 1 1170
box -8 -3 16 105
use FILL  FILL_2913
timestamp 1711653199
transform 1 0 272 0 1 1170
box -8 -3 16 105
use FILL  FILL_2914
timestamp 1711653199
transform 1 0 264 0 1 1170
box -8 -3 16 105
use FILL  FILL_2915
timestamp 1711653199
transform 1 0 256 0 1 1170
box -8 -3 16 105
use FILL  FILL_2916
timestamp 1711653199
transform 1 0 248 0 1 1170
box -8 -3 16 105
use FILL  FILL_2917
timestamp 1711653199
transform 1 0 240 0 1 1170
box -8 -3 16 105
use FILL  FILL_2918
timestamp 1711653199
transform 1 0 192 0 1 1170
box -8 -3 16 105
use FILL  FILL_2919
timestamp 1711653199
transform 1 0 184 0 1 1170
box -8 -3 16 105
use FILL  FILL_2920
timestamp 1711653199
transform 1 0 176 0 1 1170
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1711653199
transform 1 0 168 0 1 1170
box -8 -3 16 105
use FILL  FILL_2922
timestamp 1711653199
transform 1 0 160 0 1 1170
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1711653199
transform 1 0 112 0 1 1170
box -8 -3 16 105
use FILL  FILL_2924
timestamp 1711653199
transform 1 0 104 0 1 1170
box -8 -3 16 105
use FILL  FILL_2925
timestamp 1711653199
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1711653199
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1711653199
transform 1 0 3392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2928
timestamp 1711653199
transform 1 0 3384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2929
timestamp 1711653199
transform 1 0 3376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1711653199
transform 1 0 3352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2931
timestamp 1711653199
transform 1 0 3312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1711653199
transform 1 0 3304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2933
timestamp 1711653199
transform 1 0 3296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2934
timestamp 1711653199
transform 1 0 3288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1711653199
transform 1 0 3280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2936
timestamp 1711653199
transform 1 0 3272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2937
timestamp 1711653199
transform 1 0 3264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2938
timestamp 1711653199
transform 1 0 3216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2939
timestamp 1711653199
transform 1 0 3208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2940
timestamp 1711653199
transform 1 0 3200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1711653199
transform 1 0 3192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2942
timestamp 1711653199
transform 1 0 3184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1711653199
transform 1 0 3176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2944
timestamp 1711653199
transform 1 0 3168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2945
timestamp 1711653199
transform 1 0 3120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2946
timestamp 1711653199
transform 1 0 3112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2947
timestamp 1711653199
transform 1 0 3104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1711653199
transform 1 0 3096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1711653199
transform 1 0 3088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2950
timestamp 1711653199
transform 1 0 3080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2951
timestamp 1711653199
transform 1 0 3040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1711653199
transform 1 0 3032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2953
timestamp 1711653199
transform 1 0 3024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2954
timestamp 1711653199
transform 1 0 3016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2955
timestamp 1711653199
transform 1 0 2984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1711653199
transform 1 0 2976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1711653199
transform 1 0 2968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2958
timestamp 1711653199
transform 1 0 2960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2959
timestamp 1711653199
transform 1 0 2936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2960
timestamp 1711653199
transform 1 0 2928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1711653199
transform 1 0 2920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2962
timestamp 1711653199
transform 1 0 2872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1711653199
transform 1 0 2864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2964
timestamp 1711653199
transform 1 0 2856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2965
timestamp 1711653199
transform 1 0 2848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2966
timestamp 1711653199
transform 1 0 2840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2967
timestamp 1711653199
transform 1 0 2832 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2968
timestamp 1711653199
transform 1 0 2824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2969
timestamp 1711653199
transform 1 0 2768 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1711653199
transform 1 0 2760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2971
timestamp 1711653199
transform 1 0 2752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2972
timestamp 1711653199
transform 1 0 2744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2973
timestamp 1711653199
transform 1 0 2736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2974
timestamp 1711653199
transform 1 0 2728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2975
timestamp 1711653199
transform 1 0 2696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1711653199
transform 1 0 2664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2977
timestamp 1711653199
transform 1 0 2656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1711653199
transform 1 0 2648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2979
timestamp 1711653199
transform 1 0 2624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2980
timestamp 1711653199
transform 1 0 2616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2981
timestamp 1711653199
transform 1 0 2608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1711653199
transform 1 0 2568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1711653199
transform 1 0 2560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2984
timestamp 1711653199
transform 1 0 2552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1711653199
transform 1 0 2504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2986
timestamp 1711653199
transform 1 0 2496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2987
timestamp 1711653199
transform 1 0 2488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1711653199
transform 1 0 2480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2989
timestamp 1711653199
transform 1 0 2472 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2990
timestamp 1711653199
transform 1 0 2464 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1711653199
transform 1 0 2416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1711653199
transform 1 0 2408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2993
timestamp 1711653199
transform 1 0 2400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2994
timestamp 1711653199
transform 1 0 2392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2995
timestamp 1711653199
transform 1 0 2384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2996
timestamp 1711653199
transform 1 0 2376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2997
timestamp 1711653199
transform 1 0 2328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1711653199
transform 1 0 2320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1711653199
transform 1 0 2312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3000
timestamp 1711653199
transform 1 0 2304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1711653199
transform 1 0 2296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3002
timestamp 1711653199
transform 1 0 2288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3003
timestamp 1711653199
transform 1 0 2240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1711653199
transform 1 0 2232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1711653199
transform 1 0 2224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1711653199
transform 1 0 2216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1711653199
transform 1 0 2208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3008
timestamp 1711653199
transform 1 0 2176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3009
timestamp 1711653199
transform 1 0 2168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3010
timestamp 1711653199
transform 1 0 2160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1711653199
transform 1 0 2128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3012
timestamp 1711653199
transform 1 0 2120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3013
timestamp 1711653199
transform 1 0 2112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3014
timestamp 1711653199
transform 1 0 2104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3015
timestamp 1711653199
transform 1 0 2096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3016
timestamp 1711653199
transform 1 0 2048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3017
timestamp 1711653199
transform 1 0 2040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3018
timestamp 1711653199
transform 1 0 2032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3019
timestamp 1711653199
transform 1 0 2024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1711653199
transform 1 0 1984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1711653199
transform 1 0 1976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3022
timestamp 1711653199
transform 1 0 1968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3023
timestamp 1711653199
transform 1 0 1960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1711653199
transform 1 0 1952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3025
timestamp 1711653199
transform 1 0 1928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3026
timestamp 1711653199
transform 1 0 1920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3027
timestamp 1711653199
transform 1 0 1880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1711653199
transform 1 0 1872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3029
timestamp 1711653199
transform 1 0 1864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3030
timestamp 1711653199
transform 1 0 1856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1711653199
transform 1 0 1848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3032
timestamp 1711653199
transform 1 0 1824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3033
timestamp 1711653199
transform 1 0 1816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3034
timestamp 1711653199
transform 1 0 1808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1711653199
transform 1 0 1800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3036
timestamp 1711653199
transform 1 0 1792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3037
timestamp 1711653199
transform 1 0 1784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3038
timestamp 1711653199
transform 1 0 1744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3039
timestamp 1711653199
transform 1 0 1736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3040
timestamp 1711653199
transform 1 0 1728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3041
timestamp 1711653199
transform 1 0 1720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3042
timestamp 1711653199
transform 1 0 1712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3043
timestamp 1711653199
transform 1 0 1680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3044
timestamp 1711653199
transform 1 0 1672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3045
timestamp 1711653199
transform 1 0 1664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3046
timestamp 1711653199
transform 1 0 1656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1711653199
transform 1 0 1648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3048
timestamp 1711653199
transform 1 0 1640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1711653199
transform 1 0 1632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3050
timestamp 1711653199
transform 1 0 1584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3051
timestamp 1711653199
transform 1 0 1576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1711653199
transform 1 0 1568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3053
timestamp 1711653199
transform 1 0 1560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3054
timestamp 1711653199
transform 1 0 1552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3055
timestamp 1711653199
transform 1 0 1520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3056
timestamp 1711653199
transform 1 0 1512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3057
timestamp 1711653199
transform 1 0 1504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1711653199
transform 1 0 1496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3059
timestamp 1711653199
transform 1 0 1488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3060
timestamp 1711653199
transform 1 0 1480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1711653199
transform 1 0 1440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3062
timestamp 1711653199
transform 1 0 1432 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3063
timestamp 1711653199
transform 1 0 1424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3064
timestamp 1711653199
transform 1 0 1416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1711653199
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3066
timestamp 1711653199
transform 1 0 1368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1711653199
transform 1 0 1360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1711653199
transform 1 0 1352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3069
timestamp 1711653199
transform 1 0 1344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3070
timestamp 1711653199
transform 1 0 1336 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3071
timestamp 1711653199
transform 1 0 1328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1711653199
transform 1 0 1296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3073
timestamp 1711653199
transform 1 0 1288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1711653199
transform 1 0 1280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3075
timestamp 1711653199
transform 1 0 1272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3076
timestamp 1711653199
transform 1 0 1264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3077
timestamp 1711653199
transform 1 0 1216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3078
timestamp 1711653199
transform 1 0 1208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1711653199
transform 1 0 1200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3080
timestamp 1711653199
transform 1 0 1192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3081
timestamp 1711653199
transform 1 0 1184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3082
timestamp 1711653199
transform 1 0 1152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1711653199
transform 1 0 1144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3084
timestamp 1711653199
transform 1 0 1136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3085
timestamp 1711653199
transform 1 0 1128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1711653199
transform 1 0 1120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3087
timestamp 1711653199
transform 1 0 1072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3088
timestamp 1711653199
transform 1 0 1064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1711653199
transform 1 0 1056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1711653199
transform 1 0 1048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3091
timestamp 1711653199
transform 1 0 1040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3092
timestamp 1711653199
transform 1 0 1008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3093
timestamp 1711653199
transform 1 0 1000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3094
timestamp 1711653199
transform 1 0 968 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3095
timestamp 1711653199
transform 1 0 960 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3096
timestamp 1711653199
transform 1 0 952 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3097
timestamp 1711653199
transform 1 0 928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3098
timestamp 1711653199
transform 1 0 920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3099
timestamp 1711653199
transform 1 0 912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3100
timestamp 1711653199
transform 1 0 880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1711653199
transform 1 0 872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3102
timestamp 1711653199
transform 1 0 864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1711653199
transform 1 0 840 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3104
timestamp 1711653199
transform 1 0 808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3105
timestamp 1711653199
transform 1 0 800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1711653199
transform 1 0 792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3107
timestamp 1711653199
transform 1 0 760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3108
timestamp 1711653199
transform 1 0 752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3109
timestamp 1711653199
transform 1 0 744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3110
timestamp 1711653199
transform 1 0 696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1711653199
transform 1 0 688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1711653199
transform 1 0 680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3113
timestamp 1711653199
transform 1 0 672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3114
timestamp 1711653199
transform 1 0 624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3115
timestamp 1711653199
transform 1 0 616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1711653199
transform 1 0 608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3117
timestamp 1711653199
transform 1 0 600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1711653199
transform 1 0 592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3119
timestamp 1711653199
transform 1 0 544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3120
timestamp 1711653199
transform 1 0 536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1711653199
transform 1 0 504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1711653199
transform 1 0 496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3123
timestamp 1711653199
transform 1 0 488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3124
timestamp 1711653199
transform 1 0 456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3125
timestamp 1711653199
transform 1 0 448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3126
timestamp 1711653199
transform 1 0 440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1711653199
transform 1 0 392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3128
timestamp 1711653199
transform 1 0 384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3129
timestamp 1711653199
transform 1 0 376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3130
timestamp 1711653199
transform 1 0 368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3131
timestamp 1711653199
transform 1 0 320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3132
timestamp 1711653199
transform 1 0 312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3133
timestamp 1711653199
transform 1 0 280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3134
timestamp 1711653199
transform 1 0 272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3135
timestamp 1711653199
transform 1 0 264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3136
timestamp 1711653199
transform 1 0 256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3137
timestamp 1711653199
transform 1 0 248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3138
timestamp 1711653199
transform 1 0 192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3139
timestamp 1711653199
transform 1 0 184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3140
timestamp 1711653199
transform 1 0 176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3141
timestamp 1711653199
transform 1 0 136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3142
timestamp 1711653199
transform 1 0 128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3143
timestamp 1711653199
transform 1 0 88 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3144
timestamp 1711653199
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3145
timestamp 1711653199
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3146
timestamp 1711653199
transform 1 0 3392 0 1 970
box -8 -3 16 105
use FILL  FILL_3147
timestamp 1711653199
transform 1 0 3384 0 1 970
box -8 -3 16 105
use FILL  FILL_3148
timestamp 1711653199
transform 1 0 3376 0 1 970
box -8 -3 16 105
use FILL  FILL_3149
timestamp 1711653199
transform 1 0 3368 0 1 970
box -8 -3 16 105
use FILL  FILL_3150
timestamp 1711653199
transform 1 0 3360 0 1 970
box -8 -3 16 105
use FILL  FILL_3151
timestamp 1711653199
transform 1 0 3352 0 1 970
box -8 -3 16 105
use FILL  FILL_3152
timestamp 1711653199
transform 1 0 3320 0 1 970
box -8 -3 16 105
use FILL  FILL_3153
timestamp 1711653199
transform 1 0 3312 0 1 970
box -8 -3 16 105
use FILL  FILL_3154
timestamp 1711653199
transform 1 0 3304 0 1 970
box -8 -3 16 105
use FILL  FILL_3155
timestamp 1711653199
transform 1 0 3264 0 1 970
box -8 -3 16 105
use FILL  FILL_3156
timestamp 1711653199
transform 1 0 3256 0 1 970
box -8 -3 16 105
use FILL  FILL_3157
timestamp 1711653199
transform 1 0 3248 0 1 970
box -8 -3 16 105
use FILL  FILL_3158
timestamp 1711653199
transform 1 0 3240 0 1 970
box -8 -3 16 105
use FILL  FILL_3159
timestamp 1711653199
transform 1 0 3232 0 1 970
box -8 -3 16 105
use FILL  FILL_3160
timestamp 1711653199
transform 1 0 3200 0 1 970
box -8 -3 16 105
use FILL  FILL_3161
timestamp 1711653199
transform 1 0 3192 0 1 970
box -8 -3 16 105
use FILL  FILL_3162
timestamp 1711653199
transform 1 0 3184 0 1 970
box -8 -3 16 105
use FILL  FILL_3163
timestamp 1711653199
transform 1 0 3176 0 1 970
box -8 -3 16 105
use FILL  FILL_3164
timestamp 1711653199
transform 1 0 3136 0 1 970
box -8 -3 16 105
use FILL  FILL_3165
timestamp 1711653199
transform 1 0 3128 0 1 970
box -8 -3 16 105
use FILL  FILL_3166
timestamp 1711653199
transform 1 0 3120 0 1 970
box -8 -3 16 105
use FILL  FILL_3167
timestamp 1711653199
transform 1 0 3112 0 1 970
box -8 -3 16 105
use FILL  FILL_3168
timestamp 1711653199
transform 1 0 3104 0 1 970
box -8 -3 16 105
use FILL  FILL_3169
timestamp 1711653199
transform 1 0 3080 0 1 970
box -8 -3 16 105
use FILL  FILL_3170
timestamp 1711653199
transform 1 0 3072 0 1 970
box -8 -3 16 105
use FILL  FILL_3171
timestamp 1711653199
transform 1 0 3064 0 1 970
box -8 -3 16 105
use FILL  FILL_3172
timestamp 1711653199
transform 1 0 3056 0 1 970
box -8 -3 16 105
use FILL  FILL_3173
timestamp 1711653199
transform 1 0 3048 0 1 970
box -8 -3 16 105
use FILL  FILL_3174
timestamp 1711653199
transform 1 0 3008 0 1 970
box -8 -3 16 105
use FILL  FILL_3175
timestamp 1711653199
transform 1 0 3000 0 1 970
box -8 -3 16 105
use FILL  FILL_3176
timestamp 1711653199
transform 1 0 2992 0 1 970
box -8 -3 16 105
use FILL  FILL_3177
timestamp 1711653199
transform 1 0 2984 0 1 970
box -8 -3 16 105
use FILL  FILL_3178
timestamp 1711653199
transform 1 0 2976 0 1 970
box -8 -3 16 105
use FILL  FILL_3179
timestamp 1711653199
transform 1 0 2968 0 1 970
box -8 -3 16 105
use FILL  FILL_3180
timestamp 1711653199
transform 1 0 2920 0 1 970
box -8 -3 16 105
use FILL  FILL_3181
timestamp 1711653199
transform 1 0 2912 0 1 970
box -8 -3 16 105
use FILL  FILL_3182
timestamp 1711653199
transform 1 0 2904 0 1 970
box -8 -3 16 105
use FILL  FILL_3183
timestamp 1711653199
transform 1 0 2896 0 1 970
box -8 -3 16 105
use FILL  FILL_3184
timestamp 1711653199
transform 1 0 2888 0 1 970
box -8 -3 16 105
use FILL  FILL_3185
timestamp 1711653199
transform 1 0 2880 0 1 970
box -8 -3 16 105
use FILL  FILL_3186
timestamp 1711653199
transform 1 0 2840 0 1 970
box -8 -3 16 105
use FILL  FILL_3187
timestamp 1711653199
transform 1 0 2832 0 1 970
box -8 -3 16 105
use FILL  FILL_3188
timestamp 1711653199
transform 1 0 2800 0 1 970
box -8 -3 16 105
use FILL  FILL_3189
timestamp 1711653199
transform 1 0 2792 0 1 970
box -8 -3 16 105
use FILL  FILL_3190
timestamp 1711653199
transform 1 0 2784 0 1 970
box -8 -3 16 105
use FILL  FILL_3191
timestamp 1711653199
transform 1 0 2776 0 1 970
box -8 -3 16 105
use FILL  FILL_3192
timestamp 1711653199
transform 1 0 2768 0 1 970
box -8 -3 16 105
use FILL  FILL_3193
timestamp 1711653199
transform 1 0 2736 0 1 970
box -8 -3 16 105
use FILL  FILL_3194
timestamp 1711653199
transform 1 0 2728 0 1 970
box -8 -3 16 105
use FILL  FILL_3195
timestamp 1711653199
transform 1 0 2720 0 1 970
box -8 -3 16 105
use FILL  FILL_3196
timestamp 1711653199
transform 1 0 2712 0 1 970
box -8 -3 16 105
use FILL  FILL_3197
timestamp 1711653199
transform 1 0 2688 0 1 970
box -8 -3 16 105
use FILL  FILL_3198
timestamp 1711653199
transform 1 0 2656 0 1 970
box -8 -3 16 105
use FILL  FILL_3199
timestamp 1711653199
transform 1 0 2648 0 1 970
box -8 -3 16 105
use FILL  FILL_3200
timestamp 1711653199
transform 1 0 2640 0 1 970
box -8 -3 16 105
use FILL  FILL_3201
timestamp 1711653199
transform 1 0 2632 0 1 970
box -8 -3 16 105
use FILL  FILL_3202
timestamp 1711653199
transform 1 0 2624 0 1 970
box -8 -3 16 105
use FILL  FILL_3203
timestamp 1711653199
transform 1 0 2616 0 1 970
box -8 -3 16 105
use FILL  FILL_3204
timestamp 1711653199
transform 1 0 2584 0 1 970
box -8 -3 16 105
use FILL  FILL_3205
timestamp 1711653199
transform 1 0 2576 0 1 970
box -8 -3 16 105
use FILL  FILL_3206
timestamp 1711653199
transform 1 0 2544 0 1 970
box -8 -3 16 105
use FILL  FILL_3207
timestamp 1711653199
transform 1 0 2536 0 1 970
box -8 -3 16 105
use FILL  FILL_3208
timestamp 1711653199
transform 1 0 2528 0 1 970
box -8 -3 16 105
use FILL  FILL_3209
timestamp 1711653199
transform 1 0 2496 0 1 970
box -8 -3 16 105
use FILL  FILL_3210
timestamp 1711653199
transform 1 0 2488 0 1 970
box -8 -3 16 105
use FILL  FILL_3211
timestamp 1711653199
transform 1 0 2480 0 1 970
box -8 -3 16 105
use FILL  FILL_3212
timestamp 1711653199
transform 1 0 2472 0 1 970
box -8 -3 16 105
use FILL  FILL_3213
timestamp 1711653199
transform 1 0 2440 0 1 970
box -8 -3 16 105
use FILL  FILL_3214
timestamp 1711653199
transform 1 0 2432 0 1 970
box -8 -3 16 105
use FILL  FILL_3215
timestamp 1711653199
transform 1 0 2424 0 1 970
box -8 -3 16 105
use FILL  FILL_3216
timestamp 1711653199
transform 1 0 2392 0 1 970
box -8 -3 16 105
use FILL  FILL_3217
timestamp 1711653199
transform 1 0 2384 0 1 970
box -8 -3 16 105
use FILL  FILL_3218
timestamp 1711653199
transform 1 0 2376 0 1 970
box -8 -3 16 105
use FILL  FILL_3219
timestamp 1711653199
transform 1 0 2368 0 1 970
box -8 -3 16 105
use FILL  FILL_3220
timestamp 1711653199
transform 1 0 2344 0 1 970
box -8 -3 16 105
use FILL  FILL_3221
timestamp 1711653199
transform 1 0 2336 0 1 970
box -8 -3 16 105
use FILL  FILL_3222
timestamp 1711653199
transform 1 0 2328 0 1 970
box -8 -3 16 105
use FILL  FILL_3223
timestamp 1711653199
transform 1 0 2320 0 1 970
box -8 -3 16 105
use FILL  FILL_3224
timestamp 1711653199
transform 1 0 2280 0 1 970
box -8 -3 16 105
use FILL  FILL_3225
timestamp 1711653199
transform 1 0 2272 0 1 970
box -8 -3 16 105
use FILL  FILL_3226
timestamp 1711653199
transform 1 0 2264 0 1 970
box -8 -3 16 105
use FILL  FILL_3227
timestamp 1711653199
transform 1 0 2256 0 1 970
box -8 -3 16 105
use FILL  FILL_3228
timestamp 1711653199
transform 1 0 2248 0 1 970
box -8 -3 16 105
use FILL  FILL_3229
timestamp 1711653199
transform 1 0 2240 0 1 970
box -8 -3 16 105
use FILL  FILL_3230
timestamp 1711653199
transform 1 0 2192 0 1 970
box -8 -3 16 105
use FILL  FILL_3231
timestamp 1711653199
transform 1 0 2184 0 1 970
box -8 -3 16 105
use FILL  FILL_3232
timestamp 1711653199
transform 1 0 2176 0 1 970
box -8 -3 16 105
use FILL  FILL_3233
timestamp 1711653199
transform 1 0 2168 0 1 970
box -8 -3 16 105
use FILL  FILL_3234
timestamp 1711653199
transform 1 0 2160 0 1 970
box -8 -3 16 105
use FILL  FILL_3235
timestamp 1711653199
transform 1 0 2152 0 1 970
box -8 -3 16 105
use FILL  FILL_3236
timestamp 1711653199
transform 1 0 2144 0 1 970
box -8 -3 16 105
use FILL  FILL_3237
timestamp 1711653199
transform 1 0 2088 0 1 970
box -8 -3 16 105
use FILL  FILL_3238
timestamp 1711653199
transform 1 0 2080 0 1 970
box -8 -3 16 105
use FILL  FILL_3239
timestamp 1711653199
transform 1 0 2072 0 1 970
box -8 -3 16 105
use FILL  FILL_3240
timestamp 1711653199
transform 1 0 2048 0 1 970
box -8 -3 16 105
use FILL  FILL_3241
timestamp 1711653199
transform 1 0 2040 0 1 970
box -8 -3 16 105
use FILL  FILL_3242
timestamp 1711653199
transform 1 0 2032 0 1 970
box -8 -3 16 105
use FILL  FILL_3243
timestamp 1711653199
transform 1 0 1992 0 1 970
box -8 -3 16 105
use FILL  FILL_3244
timestamp 1711653199
transform 1 0 1984 0 1 970
box -8 -3 16 105
use FILL  FILL_3245
timestamp 1711653199
transform 1 0 1976 0 1 970
box -8 -3 16 105
use FILL  FILL_3246
timestamp 1711653199
transform 1 0 1952 0 1 970
box -8 -3 16 105
use FILL  FILL_3247
timestamp 1711653199
transform 1 0 1944 0 1 970
box -8 -3 16 105
use FILL  FILL_3248
timestamp 1711653199
transform 1 0 1936 0 1 970
box -8 -3 16 105
use FILL  FILL_3249
timestamp 1711653199
transform 1 0 1928 0 1 970
box -8 -3 16 105
use FILL  FILL_3250
timestamp 1711653199
transform 1 0 1888 0 1 970
box -8 -3 16 105
use FILL  FILL_3251
timestamp 1711653199
transform 1 0 1880 0 1 970
box -8 -3 16 105
use FILL  FILL_3252
timestamp 1711653199
transform 1 0 1872 0 1 970
box -8 -3 16 105
use FILL  FILL_3253
timestamp 1711653199
transform 1 0 1864 0 1 970
box -8 -3 16 105
use FILL  FILL_3254
timestamp 1711653199
transform 1 0 1824 0 1 970
box -8 -3 16 105
use FILL  FILL_3255
timestamp 1711653199
transform 1 0 1816 0 1 970
box -8 -3 16 105
use FILL  FILL_3256
timestamp 1711653199
transform 1 0 1808 0 1 970
box -8 -3 16 105
use FILL  FILL_3257
timestamp 1711653199
transform 1 0 1800 0 1 970
box -8 -3 16 105
use FILL  FILL_3258
timestamp 1711653199
transform 1 0 1792 0 1 970
box -8 -3 16 105
use FILL  FILL_3259
timestamp 1711653199
transform 1 0 1768 0 1 970
box -8 -3 16 105
use FILL  FILL_3260
timestamp 1711653199
transform 1 0 1760 0 1 970
box -8 -3 16 105
use FILL  FILL_3261
timestamp 1711653199
transform 1 0 1752 0 1 970
box -8 -3 16 105
use FILL  FILL_3262
timestamp 1711653199
transform 1 0 1720 0 1 970
box -8 -3 16 105
use FILL  FILL_3263
timestamp 1711653199
transform 1 0 1712 0 1 970
box -8 -3 16 105
use FILL  FILL_3264
timestamp 1711653199
transform 1 0 1704 0 1 970
box -8 -3 16 105
use FILL  FILL_3265
timestamp 1711653199
transform 1 0 1696 0 1 970
box -8 -3 16 105
use FILL  FILL_3266
timestamp 1711653199
transform 1 0 1688 0 1 970
box -8 -3 16 105
use FILL  FILL_3267
timestamp 1711653199
transform 1 0 1680 0 1 970
box -8 -3 16 105
use FILL  FILL_3268
timestamp 1711653199
transform 1 0 1656 0 1 970
box -8 -3 16 105
use FILL  FILL_3269
timestamp 1711653199
transform 1 0 1648 0 1 970
box -8 -3 16 105
use FILL  FILL_3270
timestamp 1711653199
transform 1 0 1616 0 1 970
box -8 -3 16 105
use FILL  FILL_3271
timestamp 1711653199
transform 1 0 1608 0 1 970
box -8 -3 16 105
use FILL  FILL_3272
timestamp 1711653199
transform 1 0 1600 0 1 970
box -8 -3 16 105
use FILL  FILL_3273
timestamp 1711653199
transform 1 0 1592 0 1 970
box -8 -3 16 105
use FILL  FILL_3274
timestamp 1711653199
transform 1 0 1584 0 1 970
box -8 -3 16 105
use FILL  FILL_3275
timestamp 1711653199
transform 1 0 1576 0 1 970
box -8 -3 16 105
use FILL  FILL_3276
timestamp 1711653199
transform 1 0 1544 0 1 970
box -8 -3 16 105
use FILL  FILL_3277
timestamp 1711653199
transform 1 0 1536 0 1 970
box -8 -3 16 105
use FILL  FILL_3278
timestamp 1711653199
transform 1 0 1528 0 1 970
box -8 -3 16 105
use FILL  FILL_3279
timestamp 1711653199
transform 1 0 1520 0 1 970
box -8 -3 16 105
use FILL  FILL_3280
timestamp 1711653199
transform 1 0 1488 0 1 970
box -8 -3 16 105
use FILL  FILL_3281
timestamp 1711653199
transform 1 0 1480 0 1 970
box -8 -3 16 105
use FILL  FILL_3282
timestamp 1711653199
transform 1 0 1472 0 1 970
box -8 -3 16 105
use FILL  FILL_3283
timestamp 1711653199
transform 1 0 1464 0 1 970
box -8 -3 16 105
use FILL  FILL_3284
timestamp 1711653199
transform 1 0 1456 0 1 970
box -8 -3 16 105
use FILL  FILL_3285
timestamp 1711653199
transform 1 0 1424 0 1 970
box -8 -3 16 105
use FILL  FILL_3286
timestamp 1711653199
transform 1 0 1416 0 1 970
box -8 -3 16 105
use FILL  FILL_3287
timestamp 1711653199
transform 1 0 1408 0 1 970
box -8 -3 16 105
use FILL  FILL_3288
timestamp 1711653199
transform 1 0 1400 0 1 970
box -8 -3 16 105
use FILL  FILL_3289
timestamp 1711653199
transform 1 0 1368 0 1 970
box -8 -3 16 105
use FILL  FILL_3290
timestamp 1711653199
transform 1 0 1360 0 1 970
box -8 -3 16 105
use FILL  FILL_3291
timestamp 1711653199
transform 1 0 1352 0 1 970
box -8 -3 16 105
use FILL  FILL_3292
timestamp 1711653199
transform 1 0 1344 0 1 970
box -8 -3 16 105
use FILL  FILL_3293
timestamp 1711653199
transform 1 0 1336 0 1 970
box -8 -3 16 105
use FILL  FILL_3294
timestamp 1711653199
transform 1 0 1328 0 1 970
box -8 -3 16 105
use FILL  FILL_3295
timestamp 1711653199
transform 1 0 1320 0 1 970
box -8 -3 16 105
use FILL  FILL_3296
timestamp 1711653199
transform 1 0 1272 0 1 970
box -8 -3 16 105
use FILL  FILL_3297
timestamp 1711653199
transform 1 0 1264 0 1 970
box -8 -3 16 105
use FILL  FILL_3298
timestamp 1711653199
transform 1 0 1256 0 1 970
box -8 -3 16 105
use FILL  FILL_3299
timestamp 1711653199
transform 1 0 1248 0 1 970
box -8 -3 16 105
use FILL  FILL_3300
timestamp 1711653199
transform 1 0 1224 0 1 970
box -8 -3 16 105
use FILL  FILL_3301
timestamp 1711653199
transform 1 0 1216 0 1 970
box -8 -3 16 105
use FILL  FILL_3302
timestamp 1711653199
transform 1 0 1208 0 1 970
box -8 -3 16 105
use FILL  FILL_3303
timestamp 1711653199
transform 1 0 1200 0 1 970
box -8 -3 16 105
use FILL  FILL_3304
timestamp 1711653199
transform 1 0 1192 0 1 970
box -8 -3 16 105
use FILL  FILL_3305
timestamp 1711653199
transform 1 0 1152 0 1 970
box -8 -3 16 105
use FILL  FILL_3306
timestamp 1711653199
transform 1 0 1144 0 1 970
box -8 -3 16 105
use FILL  FILL_3307
timestamp 1711653199
transform 1 0 1136 0 1 970
box -8 -3 16 105
use FILL  FILL_3308
timestamp 1711653199
transform 1 0 1104 0 1 970
box -8 -3 16 105
use FILL  FILL_3309
timestamp 1711653199
transform 1 0 1096 0 1 970
box -8 -3 16 105
use FILL  FILL_3310
timestamp 1711653199
transform 1 0 1088 0 1 970
box -8 -3 16 105
use FILL  FILL_3311
timestamp 1711653199
transform 1 0 1080 0 1 970
box -8 -3 16 105
use FILL  FILL_3312
timestamp 1711653199
transform 1 0 1072 0 1 970
box -8 -3 16 105
use FILL  FILL_3313
timestamp 1711653199
transform 1 0 1024 0 1 970
box -8 -3 16 105
use FILL  FILL_3314
timestamp 1711653199
transform 1 0 1016 0 1 970
box -8 -3 16 105
use FILL  FILL_3315
timestamp 1711653199
transform 1 0 1008 0 1 970
box -8 -3 16 105
use FILL  FILL_3316
timestamp 1711653199
transform 1 0 1000 0 1 970
box -8 -3 16 105
use FILL  FILL_3317
timestamp 1711653199
transform 1 0 992 0 1 970
box -8 -3 16 105
use FILL  FILL_3318
timestamp 1711653199
transform 1 0 944 0 1 970
box -8 -3 16 105
use FILL  FILL_3319
timestamp 1711653199
transform 1 0 936 0 1 970
box -8 -3 16 105
use FILL  FILL_3320
timestamp 1711653199
transform 1 0 928 0 1 970
box -8 -3 16 105
use FILL  FILL_3321
timestamp 1711653199
transform 1 0 920 0 1 970
box -8 -3 16 105
use FILL  FILL_3322
timestamp 1711653199
transform 1 0 912 0 1 970
box -8 -3 16 105
use FILL  FILL_3323
timestamp 1711653199
transform 1 0 904 0 1 970
box -8 -3 16 105
use FILL  FILL_3324
timestamp 1711653199
transform 1 0 896 0 1 970
box -8 -3 16 105
use FILL  FILL_3325
timestamp 1711653199
transform 1 0 840 0 1 970
box -8 -3 16 105
use FILL  FILL_3326
timestamp 1711653199
transform 1 0 832 0 1 970
box -8 -3 16 105
use FILL  FILL_3327
timestamp 1711653199
transform 1 0 824 0 1 970
box -8 -3 16 105
use FILL  FILL_3328
timestamp 1711653199
transform 1 0 816 0 1 970
box -8 -3 16 105
use FILL  FILL_3329
timestamp 1711653199
transform 1 0 768 0 1 970
box -8 -3 16 105
use FILL  FILL_3330
timestamp 1711653199
transform 1 0 760 0 1 970
box -8 -3 16 105
use FILL  FILL_3331
timestamp 1711653199
transform 1 0 752 0 1 970
box -8 -3 16 105
use FILL  FILL_3332
timestamp 1711653199
transform 1 0 744 0 1 970
box -8 -3 16 105
use FILL  FILL_3333
timestamp 1711653199
transform 1 0 736 0 1 970
box -8 -3 16 105
use FILL  FILL_3334
timestamp 1711653199
transform 1 0 728 0 1 970
box -8 -3 16 105
use FILL  FILL_3335
timestamp 1711653199
transform 1 0 720 0 1 970
box -8 -3 16 105
use FILL  FILL_3336
timestamp 1711653199
transform 1 0 672 0 1 970
box -8 -3 16 105
use FILL  FILL_3337
timestamp 1711653199
transform 1 0 664 0 1 970
box -8 -3 16 105
use FILL  FILL_3338
timestamp 1711653199
transform 1 0 656 0 1 970
box -8 -3 16 105
use FILL  FILL_3339
timestamp 1711653199
transform 1 0 648 0 1 970
box -8 -3 16 105
use FILL  FILL_3340
timestamp 1711653199
transform 1 0 608 0 1 970
box -8 -3 16 105
use FILL  FILL_3341
timestamp 1711653199
transform 1 0 600 0 1 970
box -8 -3 16 105
use FILL  FILL_3342
timestamp 1711653199
transform 1 0 592 0 1 970
box -8 -3 16 105
use FILL  FILL_3343
timestamp 1711653199
transform 1 0 552 0 1 970
box -8 -3 16 105
use FILL  FILL_3344
timestamp 1711653199
transform 1 0 544 0 1 970
box -8 -3 16 105
use FILL  FILL_3345
timestamp 1711653199
transform 1 0 536 0 1 970
box -8 -3 16 105
use FILL  FILL_3346
timestamp 1711653199
transform 1 0 528 0 1 970
box -8 -3 16 105
use FILL  FILL_3347
timestamp 1711653199
transform 1 0 504 0 1 970
box -8 -3 16 105
use FILL  FILL_3348
timestamp 1711653199
transform 1 0 496 0 1 970
box -8 -3 16 105
use FILL  FILL_3349
timestamp 1711653199
transform 1 0 488 0 1 970
box -8 -3 16 105
use FILL  FILL_3350
timestamp 1711653199
transform 1 0 440 0 1 970
box -8 -3 16 105
use FILL  FILL_3351
timestamp 1711653199
transform 1 0 432 0 1 970
box -8 -3 16 105
use FILL  FILL_3352
timestamp 1711653199
transform 1 0 424 0 1 970
box -8 -3 16 105
use FILL  FILL_3353
timestamp 1711653199
transform 1 0 416 0 1 970
box -8 -3 16 105
use FILL  FILL_3354
timestamp 1711653199
transform 1 0 376 0 1 970
box -8 -3 16 105
use FILL  FILL_3355
timestamp 1711653199
transform 1 0 368 0 1 970
box -8 -3 16 105
use FILL  FILL_3356
timestamp 1711653199
transform 1 0 360 0 1 970
box -8 -3 16 105
use FILL  FILL_3357
timestamp 1711653199
transform 1 0 352 0 1 970
box -8 -3 16 105
use FILL  FILL_3358
timestamp 1711653199
transform 1 0 320 0 1 970
box -8 -3 16 105
use FILL  FILL_3359
timestamp 1711653199
transform 1 0 280 0 1 970
box -8 -3 16 105
use FILL  FILL_3360
timestamp 1711653199
transform 1 0 272 0 1 970
box -8 -3 16 105
use FILL  FILL_3361
timestamp 1711653199
transform 1 0 264 0 1 970
box -8 -3 16 105
use FILL  FILL_3362
timestamp 1711653199
transform 1 0 256 0 1 970
box -8 -3 16 105
use FILL  FILL_3363
timestamp 1711653199
transform 1 0 248 0 1 970
box -8 -3 16 105
use FILL  FILL_3364
timestamp 1711653199
transform 1 0 216 0 1 970
box -8 -3 16 105
use FILL  FILL_3365
timestamp 1711653199
transform 1 0 184 0 1 970
box -8 -3 16 105
use FILL  FILL_3366
timestamp 1711653199
transform 1 0 176 0 1 970
box -8 -3 16 105
use FILL  FILL_3367
timestamp 1711653199
transform 1 0 168 0 1 970
box -8 -3 16 105
use FILL  FILL_3368
timestamp 1711653199
transform 1 0 160 0 1 970
box -8 -3 16 105
use FILL  FILL_3369
timestamp 1711653199
transform 1 0 152 0 1 970
box -8 -3 16 105
use FILL  FILL_3370
timestamp 1711653199
transform 1 0 144 0 1 970
box -8 -3 16 105
use FILL  FILL_3371
timestamp 1711653199
transform 1 0 136 0 1 970
box -8 -3 16 105
use FILL  FILL_3372
timestamp 1711653199
transform 1 0 80 0 1 970
box -8 -3 16 105
use FILL  FILL_3373
timestamp 1711653199
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_3374
timestamp 1711653199
transform 1 0 3392 0 -1 970
box -8 -3 16 105
use FILL  FILL_3375
timestamp 1711653199
transform 1 0 3384 0 -1 970
box -8 -3 16 105
use FILL  FILL_3376
timestamp 1711653199
transform 1 0 3376 0 -1 970
box -8 -3 16 105
use FILL  FILL_3377
timestamp 1711653199
transform 1 0 3320 0 -1 970
box -8 -3 16 105
use FILL  FILL_3378
timestamp 1711653199
transform 1 0 3312 0 -1 970
box -8 -3 16 105
use FILL  FILL_3379
timestamp 1711653199
transform 1 0 3304 0 -1 970
box -8 -3 16 105
use FILL  FILL_3380
timestamp 1711653199
transform 1 0 3296 0 -1 970
box -8 -3 16 105
use FILL  FILL_3381
timestamp 1711653199
transform 1 0 3288 0 -1 970
box -8 -3 16 105
use FILL  FILL_3382
timestamp 1711653199
transform 1 0 3280 0 -1 970
box -8 -3 16 105
use FILL  FILL_3383
timestamp 1711653199
transform 1 0 3232 0 -1 970
box -8 -3 16 105
use FILL  FILL_3384
timestamp 1711653199
transform 1 0 3224 0 -1 970
box -8 -3 16 105
use FILL  FILL_3385
timestamp 1711653199
transform 1 0 3216 0 -1 970
box -8 -3 16 105
use FILL  FILL_3386
timestamp 1711653199
transform 1 0 3208 0 -1 970
box -8 -3 16 105
use FILL  FILL_3387
timestamp 1711653199
transform 1 0 3176 0 -1 970
box -8 -3 16 105
use FILL  FILL_3388
timestamp 1711653199
transform 1 0 3168 0 -1 970
box -8 -3 16 105
use FILL  FILL_3389
timestamp 1711653199
transform 1 0 3160 0 -1 970
box -8 -3 16 105
use FILL  FILL_3390
timestamp 1711653199
transform 1 0 3112 0 -1 970
box -8 -3 16 105
use FILL  FILL_3391
timestamp 1711653199
transform 1 0 3104 0 -1 970
box -8 -3 16 105
use FILL  FILL_3392
timestamp 1711653199
transform 1 0 3096 0 -1 970
box -8 -3 16 105
use FILL  FILL_3393
timestamp 1711653199
transform 1 0 3088 0 -1 970
box -8 -3 16 105
use FILL  FILL_3394
timestamp 1711653199
transform 1 0 3080 0 -1 970
box -8 -3 16 105
use FILL  FILL_3395
timestamp 1711653199
transform 1 0 3072 0 -1 970
box -8 -3 16 105
use FILL  FILL_3396
timestamp 1711653199
transform 1 0 3032 0 -1 970
box -8 -3 16 105
use FILL  FILL_3397
timestamp 1711653199
transform 1 0 3024 0 -1 970
box -8 -3 16 105
use FILL  FILL_3398
timestamp 1711653199
transform 1 0 2992 0 -1 970
box -8 -3 16 105
use FILL  FILL_3399
timestamp 1711653199
transform 1 0 2984 0 -1 970
box -8 -3 16 105
use FILL  FILL_3400
timestamp 1711653199
transform 1 0 2976 0 -1 970
box -8 -3 16 105
use FILL  FILL_3401
timestamp 1711653199
transform 1 0 2968 0 -1 970
box -8 -3 16 105
use FILL  FILL_3402
timestamp 1711653199
transform 1 0 2944 0 -1 970
box -8 -3 16 105
use FILL  FILL_3403
timestamp 1711653199
transform 1 0 2936 0 -1 970
box -8 -3 16 105
use FILL  FILL_3404
timestamp 1711653199
transform 1 0 2896 0 -1 970
box -8 -3 16 105
use FILL  FILL_3405
timestamp 1711653199
transform 1 0 2888 0 -1 970
box -8 -3 16 105
use FILL  FILL_3406
timestamp 1711653199
transform 1 0 2880 0 -1 970
box -8 -3 16 105
use FILL  FILL_3407
timestamp 1711653199
transform 1 0 2872 0 -1 970
box -8 -3 16 105
use FILL  FILL_3408
timestamp 1711653199
transform 1 0 2832 0 -1 970
box -8 -3 16 105
use FILL  FILL_3409
timestamp 1711653199
transform 1 0 2824 0 -1 970
box -8 -3 16 105
use FILL  FILL_3410
timestamp 1711653199
transform 1 0 2792 0 -1 970
box -8 -3 16 105
use FILL  FILL_3411
timestamp 1711653199
transform 1 0 2784 0 -1 970
box -8 -3 16 105
use FILL  FILL_3412
timestamp 1711653199
transform 1 0 2776 0 -1 970
box -8 -3 16 105
use FILL  FILL_3413
timestamp 1711653199
transform 1 0 2768 0 -1 970
box -8 -3 16 105
use FILL  FILL_3414
timestamp 1711653199
transform 1 0 2704 0 -1 970
box -8 -3 16 105
use FILL  FILL_3415
timestamp 1711653199
transform 1 0 2696 0 -1 970
box -8 -3 16 105
use FILL  FILL_3416
timestamp 1711653199
transform 1 0 2688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3417
timestamp 1711653199
transform 1 0 2680 0 -1 970
box -8 -3 16 105
use FILL  FILL_3418
timestamp 1711653199
transform 1 0 2672 0 -1 970
box -8 -3 16 105
use FILL  FILL_3419
timestamp 1711653199
transform 1 0 2600 0 -1 970
box -8 -3 16 105
use FILL  FILL_3420
timestamp 1711653199
transform 1 0 2592 0 -1 970
box -8 -3 16 105
use FILL  FILL_3421
timestamp 1711653199
transform 1 0 2584 0 -1 970
box -8 -3 16 105
use FILL  FILL_3422
timestamp 1711653199
transform 1 0 2576 0 -1 970
box -8 -3 16 105
use FILL  FILL_3423
timestamp 1711653199
transform 1 0 2568 0 -1 970
box -8 -3 16 105
use FILL  FILL_3424
timestamp 1711653199
transform 1 0 2560 0 -1 970
box -8 -3 16 105
use FILL  FILL_3425
timestamp 1711653199
transform 1 0 2512 0 -1 970
box -8 -3 16 105
use FILL  FILL_3426
timestamp 1711653199
transform 1 0 2504 0 -1 970
box -8 -3 16 105
use FILL  FILL_3427
timestamp 1711653199
transform 1 0 2496 0 -1 970
box -8 -3 16 105
use FILL  FILL_3428
timestamp 1711653199
transform 1 0 2456 0 -1 970
box -8 -3 16 105
use FILL  FILL_3429
timestamp 1711653199
transform 1 0 2448 0 -1 970
box -8 -3 16 105
use FILL  FILL_3430
timestamp 1711653199
transform 1 0 2440 0 -1 970
box -8 -3 16 105
use FILL  FILL_3431
timestamp 1711653199
transform 1 0 2432 0 -1 970
box -8 -3 16 105
use FILL  FILL_3432
timestamp 1711653199
transform 1 0 2424 0 -1 970
box -8 -3 16 105
use FILL  FILL_3433
timestamp 1711653199
transform 1 0 2376 0 -1 970
box -8 -3 16 105
use FILL  FILL_3434
timestamp 1711653199
transform 1 0 2368 0 -1 970
box -8 -3 16 105
use FILL  FILL_3435
timestamp 1711653199
transform 1 0 2360 0 -1 970
box -8 -3 16 105
use FILL  FILL_3436
timestamp 1711653199
transform 1 0 2352 0 -1 970
box -8 -3 16 105
use FILL  FILL_3437
timestamp 1711653199
transform 1 0 2344 0 -1 970
box -8 -3 16 105
use FILL  FILL_3438
timestamp 1711653199
transform 1 0 2312 0 -1 970
box -8 -3 16 105
use FILL  FILL_3439
timestamp 1711653199
transform 1 0 2304 0 -1 970
box -8 -3 16 105
use FILL  FILL_3440
timestamp 1711653199
transform 1 0 2272 0 -1 970
box -8 -3 16 105
use FILL  FILL_3441
timestamp 1711653199
transform 1 0 2264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3442
timestamp 1711653199
transform 1 0 2256 0 -1 970
box -8 -3 16 105
use FILL  FILL_3443
timestamp 1711653199
transform 1 0 2248 0 -1 970
box -8 -3 16 105
use FILL  FILL_3444
timestamp 1711653199
transform 1 0 2240 0 -1 970
box -8 -3 16 105
use FILL  FILL_3445
timestamp 1711653199
transform 1 0 2192 0 -1 970
box -8 -3 16 105
use FILL  FILL_3446
timestamp 1711653199
transform 1 0 2184 0 -1 970
box -8 -3 16 105
use FILL  FILL_3447
timestamp 1711653199
transform 1 0 2176 0 -1 970
box -8 -3 16 105
use FILL  FILL_3448
timestamp 1711653199
transform 1 0 2168 0 -1 970
box -8 -3 16 105
use FILL  FILL_3449
timestamp 1711653199
transform 1 0 2160 0 -1 970
box -8 -3 16 105
use FILL  FILL_3450
timestamp 1711653199
transform 1 0 2120 0 -1 970
box -8 -3 16 105
use FILL  FILL_3451
timestamp 1711653199
transform 1 0 2112 0 -1 970
box -8 -3 16 105
use FILL  FILL_3452
timestamp 1711653199
transform 1 0 2104 0 -1 970
box -8 -3 16 105
use FILL  FILL_3453
timestamp 1711653199
transform 1 0 2096 0 -1 970
box -8 -3 16 105
use FILL  FILL_3454
timestamp 1711653199
transform 1 0 2088 0 -1 970
box -8 -3 16 105
use FILL  FILL_3455
timestamp 1711653199
transform 1 0 2040 0 -1 970
box -8 -3 16 105
use FILL  FILL_3456
timestamp 1711653199
transform 1 0 2032 0 -1 970
box -8 -3 16 105
use FILL  FILL_3457
timestamp 1711653199
transform 1 0 2024 0 -1 970
box -8 -3 16 105
use FILL  FILL_3458
timestamp 1711653199
transform 1 0 1984 0 -1 970
box -8 -3 16 105
use FILL  FILL_3459
timestamp 1711653199
transform 1 0 1976 0 -1 970
box -8 -3 16 105
use FILL  FILL_3460
timestamp 1711653199
transform 1 0 1968 0 -1 970
box -8 -3 16 105
use FILL  FILL_3461
timestamp 1711653199
transform 1 0 1928 0 -1 970
box -8 -3 16 105
use FILL  FILL_3462
timestamp 1711653199
transform 1 0 1920 0 -1 970
box -8 -3 16 105
use FILL  FILL_3463
timestamp 1711653199
transform 1 0 1912 0 -1 970
box -8 -3 16 105
use FILL  FILL_3464
timestamp 1711653199
transform 1 0 1872 0 -1 970
box -8 -3 16 105
use FILL  FILL_3465
timestamp 1711653199
transform 1 0 1864 0 -1 970
box -8 -3 16 105
use FILL  FILL_3466
timestamp 1711653199
transform 1 0 1856 0 -1 970
box -8 -3 16 105
use FILL  FILL_3467
timestamp 1711653199
transform 1 0 1848 0 -1 970
box -8 -3 16 105
use FILL  FILL_3468
timestamp 1711653199
transform 1 0 1824 0 -1 970
box -8 -3 16 105
use FILL  FILL_3469
timestamp 1711653199
transform 1 0 1784 0 -1 970
box -8 -3 16 105
use FILL  FILL_3470
timestamp 1711653199
transform 1 0 1776 0 -1 970
box -8 -3 16 105
use FILL  FILL_3471
timestamp 1711653199
transform 1 0 1768 0 -1 970
box -8 -3 16 105
use FILL  FILL_3472
timestamp 1711653199
transform 1 0 1760 0 -1 970
box -8 -3 16 105
use FILL  FILL_3473
timestamp 1711653199
transform 1 0 1752 0 -1 970
box -8 -3 16 105
use FILL  FILL_3474
timestamp 1711653199
transform 1 0 1744 0 -1 970
box -8 -3 16 105
use FILL  FILL_3475
timestamp 1711653199
transform 1 0 1736 0 -1 970
box -8 -3 16 105
use FILL  FILL_3476
timestamp 1711653199
transform 1 0 1704 0 -1 970
box -8 -3 16 105
use FILL  FILL_3477
timestamp 1711653199
transform 1 0 1696 0 -1 970
box -8 -3 16 105
use FILL  FILL_3478
timestamp 1711653199
transform 1 0 1688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3479
timestamp 1711653199
transform 1 0 1680 0 -1 970
box -8 -3 16 105
use FILL  FILL_3480
timestamp 1711653199
transform 1 0 1648 0 -1 970
box -8 -3 16 105
use FILL  FILL_3481
timestamp 1711653199
transform 1 0 1640 0 -1 970
box -8 -3 16 105
use FILL  FILL_3482
timestamp 1711653199
transform 1 0 1632 0 -1 970
box -8 -3 16 105
use FILL  FILL_3483
timestamp 1711653199
transform 1 0 1624 0 -1 970
box -8 -3 16 105
use FILL  FILL_3484
timestamp 1711653199
transform 1 0 1616 0 -1 970
box -8 -3 16 105
use FILL  FILL_3485
timestamp 1711653199
transform 1 0 1584 0 -1 970
box -8 -3 16 105
use FILL  FILL_3486
timestamp 1711653199
transform 1 0 1576 0 -1 970
box -8 -3 16 105
use FILL  FILL_3487
timestamp 1711653199
transform 1 0 1568 0 -1 970
box -8 -3 16 105
use FILL  FILL_3488
timestamp 1711653199
transform 1 0 1560 0 -1 970
box -8 -3 16 105
use FILL  FILL_3489
timestamp 1711653199
transform 1 0 1528 0 -1 970
box -8 -3 16 105
use FILL  FILL_3490
timestamp 1711653199
transform 1 0 1520 0 -1 970
box -8 -3 16 105
use FILL  FILL_3491
timestamp 1711653199
transform 1 0 1512 0 -1 970
box -8 -3 16 105
use FILL  FILL_3492
timestamp 1711653199
transform 1 0 1504 0 -1 970
box -8 -3 16 105
use FILL  FILL_3493
timestamp 1711653199
transform 1 0 1496 0 -1 970
box -8 -3 16 105
use FILL  FILL_3494
timestamp 1711653199
transform 1 0 1464 0 -1 970
box -8 -3 16 105
use FILL  FILL_3495
timestamp 1711653199
transform 1 0 1456 0 -1 970
box -8 -3 16 105
use FILL  FILL_3496
timestamp 1711653199
transform 1 0 1448 0 -1 970
box -8 -3 16 105
use FILL  FILL_3497
timestamp 1711653199
transform 1 0 1416 0 -1 970
box -8 -3 16 105
use FILL  FILL_3498
timestamp 1711653199
transform 1 0 1408 0 -1 970
box -8 -3 16 105
use FILL  FILL_3499
timestamp 1711653199
transform 1 0 1400 0 -1 970
box -8 -3 16 105
use FILL  FILL_3500
timestamp 1711653199
transform 1 0 1392 0 -1 970
box -8 -3 16 105
use FILL  FILL_3501
timestamp 1711653199
transform 1 0 1384 0 -1 970
box -8 -3 16 105
use FILL  FILL_3502
timestamp 1711653199
transform 1 0 1376 0 -1 970
box -8 -3 16 105
use FILL  FILL_3503
timestamp 1711653199
transform 1 0 1368 0 -1 970
box -8 -3 16 105
use FILL  FILL_3504
timestamp 1711653199
transform 1 0 1328 0 -1 970
box -8 -3 16 105
use FILL  FILL_3505
timestamp 1711653199
transform 1 0 1304 0 -1 970
box -8 -3 16 105
use FILL  FILL_3506
timestamp 1711653199
transform 1 0 1296 0 -1 970
box -8 -3 16 105
use FILL  FILL_3507
timestamp 1711653199
transform 1 0 1288 0 -1 970
box -8 -3 16 105
use FILL  FILL_3508
timestamp 1711653199
transform 1 0 1280 0 -1 970
box -8 -3 16 105
use FILL  FILL_3509
timestamp 1711653199
transform 1 0 1272 0 -1 970
box -8 -3 16 105
use FILL  FILL_3510
timestamp 1711653199
transform 1 0 1264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3511
timestamp 1711653199
transform 1 0 1256 0 -1 970
box -8 -3 16 105
use FILL  FILL_3512
timestamp 1711653199
transform 1 0 1208 0 -1 970
box -8 -3 16 105
use FILL  FILL_3513
timestamp 1711653199
transform 1 0 1200 0 -1 970
box -8 -3 16 105
use FILL  FILL_3514
timestamp 1711653199
transform 1 0 1192 0 -1 970
box -8 -3 16 105
use FILL  FILL_3515
timestamp 1711653199
transform 1 0 1152 0 -1 970
box -8 -3 16 105
use FILL  FILL_3516
timestamp 1711653199
transform 1 0 1144 0 -1 970
box -8 -3 16 105
use FILL  FILL_3517
timestamp 1711653199
transform 1 0 1136 0 -1 970
box -8 -3 16 105
use FILL  FILL_3518
timestamp 1711653199
transform 1 0 1128 0 -1 970
box -8 -3 16 105
use FILL  FILL_3519
timestamp 1711653199
transform 1 0 1120 0 -1 970
box -8 -3 16 105
use FILL  FILL_3520
timestamp 1711653199
transform 1 0 1072 0 -1 970
box -8 -3 16 105
use FILL  FILL_3521
timestamp 1711653199
transform 1 0 1064 0 -1 970
box -8 -3 16 105
use FILL  FILL_3522
timestamp 1711653199
transform 1 0 1056 0 -1 970
box -8 -3 16 105
use FILL  FILL_3523
timestamp 1711653199
transform 1 0 1048 0 -1 970
box -8 -3 16 105
use FILL  FILL_3524
timestamp 1711653199
transform 1 0 1024 0 -1 970
box -8 -3 16 105
use FILL  FILL_3525
timestamp 1711653199
transform 1 0 1016 0 -1 970
box -8 -3 16 105
use FILL  FILL_3526
timestamp 1711653199
transform 1 0 1008 0 -1 970
box -8 -3 16 105
use FILL  FILL_3527
timestamp 1711653199
transform 1 0 968 0 -1 970
box -8 -3 16 105
use FILL  FILL_3528
timestamp 1711653199
transform 1 0 960 0 -1 970
box -8 -3 16 105
use FILL  FILL_3529
timestamp 1711653199
transform 1 0 952 0 -1 970
box -8 -3 16 105
use FILL  FILL_3530
timestamp 1711653199
transform 1 0 944 0 -1 970
box -8 -3 16 105
use FILL  FILL_3531
timestamp 1711653199
transform 1 0 936 0 -1 970
box -8 -3 16 105
use FILL  FILL_3532
timestamp 1711653199
transform 1 0 904 0 -1 970
box -8 -3 16 105
use FILL  FILL_3533
timestamp 1711653199
transform 1 0 896 0 -1 970
box -8 -3 16 105
use FILL  FILL_3534
timestamp 1711653199
transform 1 0 872 0 -1 970
box -8 -3 16 105
use FILL  FILL_3535
timestamp 1711653199
transform 1 0 864 0 -1 970
box -8 -3 16 105
use FILL  FILL_3536
timestamp 1711653199
transform 1 0 856 0 -1 970
box -8 -3 16 105
use FILL  FILL_3537
timestamp 1711653199
transform 1 0 848 0 -1 970
box -8 -3 16 105
use FILL  FILL_3538
timestamp 1711653199
transform 1 0 824 0 -1 970
box -8 -3 16 105
use FILL  FILL_3539
timestamp 1711653199
transform 1 0 792 0 -1 970
box -8 -3 16 105
use FILL  FILL_3540
timestamp 1711653199
transform 1 0 784 0 -1 970
box -8 -3 16 105
use FILL  FILL_3541
timestamp 1711653199
transform 1 0 776 0 -1 970
box -8 -3 16 105
use FILL  FILL_3542
timestamp 1711653199
transform 1 0 768 0 -1 970
box -8 -3 16 105
use FILL  FILL_3543
timestamp 1711653199
transform 1 0 728 0 -1 970
box -8 -3 16 105
use FILL  FILL_3544
timestamp 1711653199
transform 1 0 720 0 -1 970
box -8 -3 16 105
use FILL  FILL_3545
timestamp 1711653199
transform 1 0 688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3546
timestamp 1711653199
transform 1 0 680 0 -1 970
box -8 -3 16 105
use FILL  FILL_3547
timestamp 1711653199
transform 1 0 672 0 -1 970
box -8 -3 16 105
use FILL  FILL_3548
timestamp 1711653199
transform 1 0 632 0 -1 970
box -8 -3 16 105
use FILL  FILL_3549
timestamp 1711653199
transform 1 0 624 0 -1 970
box -8 -3 16 105
use FILL  FILL_3550
timestamp 1711653199
transform 1 0 616 0 -1 970
box -8 -3 16 105
use FILL  FILL_3551
timestamp 1711653199
transform 1 0 576 0 -1 970
box -8 -3 16 105
use FILL  FILL_3552
timestamp 1711653199
transform 1 0 568 0 -1 970
box -8 -3 16 105
use FILL  FILL_3553
timestamp 1711653199
transform 1 0 560 0 -1 970
box -8 -3 16 105
use FILL  FILL_3554
timestamp 1711653199
transform 1 0 552 0 -1 970
box -8 -3 16 105
use FILL  FILL_3555
timestamp 1711653199
transform 1 0 544 0 -1 970
box -8 -3 16 105
use FILL  FILL_3556
timestamp 1711653199
transform 1 0 488 0 -1 970
box -8 -3 16 105
use FILL  FILL_3557
timestamp 1711653199
transform 1 0 480 0 -1 970
box -8 -3 16 105
use FILL  FILL_3558
timestamp 1711653199
transform 1 0 472 0 -1 970
box -8 -3 16 105
use FILL  FILL_3559
timestamp 1711653199
transform 1 0 464 0 -1 970
box -8 -3 16 105
use FILL  FILL_3560
timestamp 1711653199
transform 1 0 456 0 -1 970
box -8 -3 16 105
use FILL  FILL_3561
timestamp 1711653199
transform 1 0 416 0 -1 970
box -8 -3 16 105
use FILL  FILL_3562
timestamp 1711653199
transform 1 0 408 0 -1 970
box -8 -3 16 105
use FILL  FILL_3563
timestamp 1711653199
transform 1 0 376 0 -1 970
box -8 -3 16 105
use FILL  FILL_3564
timestamp 1711653199
transform 1 0 368 0 -1 970
box -8 -3 16 105
use FILL  FILL_3565
timestamp 1711653199
transform 1 0 360 0 -1 970
box -8 -3 16 105
use FILL  FILL_3566
timestamp 1711653199
transform 1 0 352 0 -1 970
box -8 -3 16 105
use FILL  FILL_3567
timestamp 1711653199
transform 1 0 344 0 -1 970
box -8 -3 16 105
use FILL  FILL_3568
timestamp 1711653199
transform 1 0 288 0 -1 970
box -8 -3 16 105
use FILL  FILL_3569
timestamp 1711653199
transform 1 0 280 0 -1 970
box -8 -3 16 105
use FILL  FILL_3570
timestamp 1711653199
transform 1 0 272 0 -1 970
box -8 -3 16 105
use FILL  FILL_3571
timestamp 1711653199
transform 1 0 264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3572
timestamp 1711653199
transform 1 0 256 0 -1 970
box -8 -3 16 105
use FILL  FILL_3573
timestamp 1711653199
transform 1 0 192 0 -1 970
box -8 -3 16 105
use FILL  FILL_3574
timestamp 1711653199
transform 1 0 184 0 -1 970
box -8 -3 16 105
use FILL  FILL_3575
timestamp 1711653199
transform 1 0 176 0 -1 970
box -8 -3 16 105
use FILL  FILL_3576
timestamp 1711653199
transform 1 0 168 0 -1 970
box -8 -3 16 105
use FILL  FILL_3577
timestamp 1711653199
transform 1 0 160 0 -1 970
box -8 -3 16 105
use FILL  FILL_3578
timestamp 1711653199
transform 1 0 128 0 -1 970
box -8 -3 16 105
use FILL  FILL_3579
timestamp 1711653199
transform 1 0 88 0 -1 970
box -8 -3 16 105
use FILL  FILL_3580
timestamp 1711653199
transform 1 0 80 0 -1 970
box -8 -3 16 105
use FILL  FILL_3581
timestamp 1711653199
transform 1 0 72 0 -1 970
box -8 -3 16 105
use FILL  FILL_3582
timestamp 1711653199
transform 1 0 3392 0 1 770
box -8 -3 16 105
use FILL  FILL_3583
timestamp 1711653199
transform 1 0 3384 0 1 770
box -8 -3 16 105
use FILL  FILL_3584
timestamp 1711653199
transform 1 0 3328 0 1 770
box -8 -3 16 105
use FILL  FILL_3585
timestamp 1711653199
transform 1 0 3320 0 1 770
box -8 -3 16 105
use FILL  FILL_3586
timestamp 1711653199
transform 1 0 3312 0 1 770
box -8 -3 16 105
use FILL  FILL_3587
timestamp 1711653199
transform 1 0 3304 0 1 770
box -8 -3 16 105
use FILL  FILL_3588
timestamp 1711653199
transform 1 0 3256 0 1 770
box -8 -3 16 105
use FILL  FILL_3589
timestamp 1711653199
transform 1 0 3248 0 1 770
box -8 -3 16 105
use FILL  FILL_3590
timestamp 1711653199
transform 1 0 3240 0 1 770
box -8 -3 16 105
use FILL  FILL_3591
timestamp 1711653199
transform 1 0 3192 0 1 770
box -8 -3 16 105
use FILL  FILL_3592
timestamp 1711653199
transform 1 0 3184 0 1 770
box -8 -3 16 105
use FILL  FILL_3593
timestamp 1711653199
transform 1 0 3176 0 1 770
box -8 -3 16 105
use FILL  FILL_3594
timestamp 1711653199
transform 1 0 3168 0 1 770
box -8 -3 16 105
use FILL  FILL_3595
timestamp 1711653199
transform 1 0 3160 0 1 770
box -8 -3 16 105
use FILL  FILL_3596
timestamp 1711653199
transform 1 0 3112 0 1 770
box -8 -3 16 105
use FILL  FILL_3597
timestamp 1711653199
transform 1 0 3104 0 1 770
box -8 -3 16 105
use FILL  FILL_3598
timestamp 1711653199
transform 1 0 3096 0 1 770
box -8 -3 16 105
use FILL  FILL_3599
timestamp 1711653199
transform 1 0 3088 0 1 770
box -8 -3 16 105
use FILL  FILL_3600
timestamp 1711653199
transform 1 0 3048 0 1 770
box -8 -3 16 105
use FILL  FILL_3601
timestamp 1711653199
transform 1 0 3040 0 1 770
box -8 -3 16 105
use FILL  FILL_3602
timestamp 1711653199
transform 1 0 3032 0 1 770
box -8 -3 16 105
use FILL  FILL_3603
timestamp 1711653199
transform 1 0 2992 0 1 770
box -8 -3 16 105
use FILL  FILL_3604
timestamp 1711653199
transform 1 0 2968 0 1 770
box -8 -3 16 105
use FILL  FILL_3605
timestamp 1711653199
transform 1 0 2960 0 1 770
box -8 -3 16 105
use FILL  FILL_3606
timestamp 1711653199
transform 1 0 2952 0 1 770
box -8 -3 16 105
use FILL  FILL_3607
timestamp 1711653199
transform 1 0 2944 0 1 770
box -8 -3 16 105
use FILL  FILL_3608
timestamp 1711653199
transform 1 0 2904 0 1 770
box -8 -3 16 105
use FILL  FILL_3609
timestamp 1711653199
transform 1 0 2896 0 1 770
box -8 -3 16 105
use FILL  FILL_3610
timestamp 1711653199
transform 1 0 2888 0 1 770
box -8 -3 16 105
use FILL  FILL_3611
timestamp 1711653199
transform 1 0 2848 0 1 770
box -8 -3 16 105
use FILL  FILL_3612
timestamp 1711653199
transform 1 0 2840 0 1 770
box -8 -3 16 105
use FILL  FILL_3613
timestamp 1711653199
transform 1 0 2800 0 1 770
box -8 -3 16 105
use FILL  FILL_3614
timestamp 1711653199
transform 1 0 2792 0 1 770
box -8 -3 16 105
use FILL  FILL_3615
timestamp 1711653199
transform 1 0 2784 0 1 770
box -8 -3 16 105
use FILL  FILL_3616
timestamp 1711653199
transform 1 0 2776 0 1 770
box -8 -3 16 105
use FILL  FILL_3617
timestamp 1711653199
transform 1 0 2736 0 1 770
box -8 -3 16 105
use FILL  FILL_3618
timestamp 1711653199
transform 1 0 2728 0 1 770
box -8 -3 16 105
use FILL  FILL_3619
timestamp 1711653199
transform 1 0 2720 0 1 770
box -8 -3 16 105
use FILL  FILL_3620
timestamp 1711653199
transform 1 0 2680 0 1 770
box -8 -3 16 105
use FILL  FILL_3621
timestamp 1711653199
transform 1 0 2648 0 1 770
box -8 -3 16 105
use FILL  FILL_3622
timestamp 1711653199
transform 1 0 2640 0 1 770
box -8 -3 16 105
use FILL  FILL_3623
timestamp 1711653199
transform 1 0 2632 0 1 770
box -8 -3 16 105
use FILL  FILL_3624
timestamp 1711653199
transform 1 0 2624 0 1 770
box -8 -3 16 105
use FILL  FILL_3625
timestamp 1711653199
transform 1 0 2616 0 1 770
box -8 -3 16 105
use FILL  FILL_3626
timestamp 1711653199
transform 1 0 2568 0 1 770
box -8 -3 16 105
use FILL  FILL_3627
timestamp 1711653199
transform 1 0 2560 0 1 770
box -8 -3 16 105
use FILL  FILL_3628
timestamp 1711653199
transform 1 0 2528 0 1 770
box -8 -3 16 105
use FILL  FILL_3629
timestamp 1711653199
transform 1 0 2520 0 1 770
box -8 -3 16 105
use FILL  FILL_3630
timestamp 1711653199
transform 1 0 2512 0 1 770
box -8 -3 16 105
use FILL  FILL_3631
timestamp 1711653199
transform 1 0 2504 0 1 770
box -8 -3 16 105
use FILL  FILL_3632
timestamp 1711653199
transform 1 0 2472 0 1 770
box -8 -3 16 105
use FILL  FILL_3633
timestamp 1711653199
transform 1 0 2464 0 1 770
box -8 -3 16 105
use FILL  FILL_3634
timestamp 1711653199
transform 1 0 2456 0 1 770
box -8 -3 16 105
use FILL  FILL_3635
timestamp 1711653199
transform 1 0 2408 0 1 770
box -8 -3 16 105
use FILL  FILL_3636
timestamp 1711653199
transform 1 0 2400 0 1 770
box -8 -3 16 105
use FILL  FILL_3637
timestamp 1711653199
transform 1 0 2392 0 1 770
box -8 -3 16 105
use FILL  FILL_3638
timestamp 1711653199
transform 1 0 2384 0 1 770
box -8 -3 16 105
use FILL  FILL_3639
timestamp 1711653199
transform 1 0 2376 0 1 770
box -8 -3 16 105
use FILL  FILL_3640
timestamp 1711653199
transform 1 0 2368 0 1 770
box -8 -3 16 105
use FILL  FILL_3641
timestamp 1711653199
transform 1 0 2304 0 1 770
box -8 -3 16 105
use FILL  FILL_3642
timestamp 1711653199
transform 1 0 2296 0 1 770
box -8 -3 16 105
use FILL  FILL_3643
timestamp 1711653199
transform 1 0 2288 0 1 770
box -8 -3 16 105
use FILL  FILL_3644
timestamp 1711653199
transform 1 0 2280 0 1 770
box -8 -3 16 105
use FILL  FILL_3645
timestamp 1711653199
transform 1 0 2272 0 1 770
box -8 -3 16 105
use FILL  FILL_3646
timestamp 1711653199
transform 1 0 2264 0 1 770
box -8 -3 16 105
use FILL  FILL_3647
timestamp 1711653199
transform 1 0 2232 0 1 770
box -8 -3 16 105
use FILL  FILL_3648
timestamp 1711653199
transform 1 0 2192 0 1 770
box -8 -3 16 105
use FILL  FILL_3649
timestamp 1711653199
transform 1 0 2184 0 1 770
box -8 -3 16 105
use FILL  FILL_3650
timestamp 1711653199
transform 1 0 2176 0 1 770
box -8 -3 16 105
use FILL  FILL_3651
timestamp 1711653199
transform 1 0 2168 0 1 770
box -8 -3 16 105
use FILL  FILL_3652
timestamp 1711653199
transform 1 0 2160 0 1 770
box -8 -3 16 105
use FILL  FILL_3653
timestamp 1711653199
transform 1 0 2152 0 1 770
box -8 -3 16 105
use FILL  FILL_3654
timestamp 1711653199
transform 1 0 2088 0 1 770
box -8 -3 16 105
use FILL  FILL_3655
timestamp 1711653199
transform 1 0 2080 0 1 770
box -8 -3 16 105
use FILL  FILL_3656
timestamp 1711653199
transform 1 0 2072 0 1 770
box -8 -3 16 105
use FILL  FILL_3657
timestamp 1711653199
transform 1 0 2064 0 1 770
box -8 -3 16 105
use FILL  FILL_3658
timestamp 1711653199
transform 1 0 2056 0 1 770
box -8 -3 16 105
use FILL  FILL_3659
timestamp 1711653199
transform 1 0 2000 0 1 770
box -8 -3 16 105
use FILL  FILL_3660
timestamp 1711653199
transform 1 0 1992 0 1 770
box -8 -3 16 105
use FILL  FILL_3661
timestamp 1711653199
transform 1 0 1984 0 1 770
box -8 -3 16 105
use FILL  FILL_3662
timestamp 1711653199
transform 1 0 1976 0 1 770
box -8 -3 16 105
use FILL  FILL_3663
timestamp 1711653199
transform 1 0 1928 0 1 770
box -8 -3 16 105
use FILL  FILL_3664
timestamp 1711653199
transform 1 0 1920 0 1 770
box -8 -3 16 105
use FILL  FILL_3665
timestamp 1711653199
transform 1 0 1912 0 1 770
box -8 -3 16 105
use FILL  FILL_3666
timestamp 1711653199
transform 1 0 1904 0 1 770
box -8 -3 16 105
use FILL  FILL_3667
timestamp 1711653199
transform 1 0 1896 0 1 770
box -8 -3 16 105
use FILL  FILL_3668
timestamp 1711653199
transform 1 0 1848 0 1 770
box -8 -3 16 105
use FILL  FILL_3669
timestamp 1711653199
transform 1 0 1840 0 1 770
box -8 -3 16 105
use FILL  FILL_3670
timestamp 1711653199
transform 1 0 1832 0 1 770
box -8 -3 16 105
use FILL  FILL_3671
timestamp 1711653199
transform 1 0 1824 0 1 770
box -8 -3 16 105
use FILL  FILL_3672
timestamp 1711653199
transform 1 0 1784 0 1 770
box -8 -3 16 105
use FILL  FILL_3673
timestamp 1711653199
transform 1 0 1776 0 1 770
box -8 -3 16 105
use FILL  FILL_3674
timestamp 1711653199
transform 1 0 1768 0 1 770
box -8 -3 16 105
use FILL  FILL_3675
timestamp 1711653199
transform 1 0 1760 0 1 770
box -8 -3 16 105
use FILL  FILL_3676
timestamp 1711653199
transform 1 0 1728 0 1 770
box -8 -3 16 105
use FILL  FILL_3677
timestamp 1711653199
transform 1 0 1720 0 1 770
box -8 -3 16 105
use FILL  FILL_3678
timestamp 1711653199
transform 1 0 1712 0 1 770
box -8 -3 16 105
use FILL  FILL_3679
timestamp 1711653199
transform 1 0 1680 0 1 770
box -8 -3 16 105
use FILL  FILL_3680
timestamp 1711653199
transform 1 0 1672 0 1 770
box -8 -3 16 105
use FILL  FILL_3681
timestamp 1711653199
transform 1 0 1664 0 1 770
box -8 -3 16 105
use FILL  FILL_3682
timestamp 1711653199
transform 1 0 1656 0 1 770
box -8 -3 16 105
use FILL  FILL_3683
timestamp 1711653199
transform 1 0 1608 0 1 770
box -8 -3 16 105
use FILL  FILL_3684
timestamp 1711653199
transform 1 0 1600 0 1 770
box -8 -3 16 105
use FILL  FILL_3685
timestamp 1711653199
transform 1 0 1592 0 1 770
box -8 -3 16 105
use FILL  FILL_3686
timestamp 1711653199
transform 1 0 1584 0 1 770
box -8 -3 16 105
use FILL  FILL_3687
timestamp 1711653199
transform 1 0 1576 0 1 770
box -8 -3 16 105
use FILL  FILL_3688
timestamp 1711653199
transform 1 0 1568 0 1 770
box -8 -3 16 105
use FILL  FILL_3689
timestamp 1711653199
transform 1 0 1520 0 1 770
box -8 -3 16 105
use FILL  FILL_3690
timestamp 1711653199
transform 1 0 1512 0 1 770
box -8 -3 16 105
use FILL  FILL_3691
timestamp 1711653199
transform 1 0 1504 0 1 770
box -8 -3 16 105
use FILL  FILL_3692
timestamp 1711653199
transform 1 0 1472 0 1 770
box -8 -3 16 105
use FILL  FILL_3693
timestamp 1711653199
transform 1 0 1464 0 1 770
box -8 -3 16 105
use FILL  FILL_3694
timestamp 1711653199
transform 1 0 1456 0 1 770
box -8 -3 16 105
use FILL  FILL_3695
timestamp 1711653199
transform 1 0 1448 0 1 770
box -8 -3 16 105
use FILL  FILL_3696
timestamp 1711653199
transform 1 0 1440 0 1 770
box -8 -3 16 105
use FILL  FILL_3697
timestamp 1711653199
transform 1 0 1432 0 1 770
box -8 -3 16 105
use FILL  FILL_3698
timestamp 1711653199
transform 1 0 1384 0 1 770
box -8 -3 16 105
use FILL  FILL_3699
timestamp 1711653199
transform 1 0 1376 0 1 770
box -8 -3 16 105
use FILL  FILL_3700
timestamp 1711653199
transform 1 0 1368 0 1 770
box -8 -3 16 105
use FILL  FILL_3701
timestamp 1711653199
transform 1 0 1360 0 1 770
box -8 -3 16 105
use FILL  FILL_3702
timestamp 1711653199
transform 1 0 1328 0 1 770
box -8 -3 16 105
use FILL  FILL_3703
timestamp 1711653199
transform 1 0 1320 0 1 770
box -8 -3 16 105
use FILL  FILL_3704
timestamp 1711653199
transform 1 0 1312 0 1 770
box -8 -3 16 105
use FILL  FILL_3705
timestamp 1711653199
transform 1 0 1304 0 1 770
box -8 -3 16 105
use FILL  FILL_3706
timestamp 1711653199
transform 1 0 1256 0 1 770
box -8 -3 16 105
use FILL  FILL_3707
timestamp 1711653199
transform 1 0 1248 0 1 770
box -8 -3 16 105
use FILL  FILL_3708
timestamp 1711653199
transform 1 0 1240 0 1 770
box -8 -3 16 105
use FILL  FILL_3709
timestamp 1711653199
transform 1 0 1232 0 1 770
box -8 -3 16 105
use FILL  FILL_3710
timestamp 1711653199
transform 1 0 1224 0 1 770
box -8 -3 16 105
use FILL  FILL_3711
timestamp 1711653199
transform 1 0 1216 0 1 770
box -8 -3 16 105
use FILL  FILL_3712
timestamp 1711653199
transform 1 0 1208 0 1 770
box -8 -3 16 105
use FILL  FILL_3713
timestamp 1711653199
transform 1 0 1168 0 1 770
box -8 -3 16 105
use FILL  FILL_3714
timestamp 1711653199
transform 1 0 1160 0 1 770
box -8 -3 16 105
use FILL  FILL_3715
timestamp 1711653199
transform 1 0 1152 0 1 770
box -8 -3 16 105
use FILL  FILL_3716
timestamp 1711653199
transform 1 0 1120 0 1 770
box -8 -3 16 105
use FILL  FILL_3717
timestamp 1711653199
transform 1 0 1112 0 1 770
box -8 -3 16 105
use FILL  FILL_3718
timestamp 1711653199
transform 1 0 1104 0 1 770
box -8 -3 16 105
use FILL  FILL_3719
timestamp 1711653199
transform 1 0 1096 0 1 770
box -8 -3 16 105
use FILL  FILL_3720
timestamp 1711653199
transform 1 0 1056 0 1 770
box -8 -3 16 105
use FILL  FILL_3721
timestamp 1711653199
transform 1 0 1048 0 1 770
box -8 -3 16 105
use FILL  FILL_3722
timestamp 1711653199
transform 1 0 1040 0 1 770
box -8 -3 16 105
use FILL  FILL_3723
timestamp 1711653199
transform 1 0 1032 0 1 770
box -8 -3 16 105
use FILL  FILL_3724
timestamp 1711653199
transform 1 0 1024 0 1 770
box -8 -3 16 105
use FILL  FILL_3725
timestamp 1711653199
transform 1 0 984 0 1 770
box -8 -3 16 105
use FILL  FILL_3726
timestamp 1711653199
transform 1 0 976 0 1 770
box -8 -3 16 105
use FILL  FILL_3727
timestamp 1711653199
transform 1 0 968 0 1 770
box -8 -3 16 105
use FILL  FILL_3728
timestamp 1711653199
transform 1 0 960 0 1 770
box -8 -3 16 105
use FILL  FILL_3729
timestamp 1711653199
transform 1 0 952 0 1 770
box -8 -3 16 105
use FILL  FILL_3730
timestamp 1711653199
transform 1 0 904 0 1 770
box -8 -3 16 105
use FILL  FILL_3731
timestamp 1711653199
transform 1 0 896 0 1 770
box -8 -3 16 105
use FILL  FILL_3732
timestamp 1711653199
transform 1 0 888 0 1 770
box -8 -3 16 105
use FILL  FILL_3733
timestamp 1711653199
transform 1 0 880 0 1 770
box -8 -3 16 105
use FILL  FILL_3734
timestamp 1711653199
transform 1 0 872 0 1 770
box -8 -3 16 105
use FILL  FILL_3735
timestamp 1711653199
transform 1 0 840 0 1 770
box -8 -3 16 105
use FILL  FILL_3736
timestamp 1711653199
transform 1 0 832 0 1 770
box -8 -3 16 105
use FILL  FILL_3737
timestamp 1711653199
transform 1 0 824 0 1 770
box -8 -3 16 105
use FILL  FILL_3738
timestamp 1711653199
transform 1 0 784 0 1 770
box -8 -3 16 105
use FILL  FILL_3739
timestamp 1711653199
transform 1 0 776 0 1 770
box -8 -3 16 105
use FILL  FILL_3740
timestamp 1711653199
transform 1 0 768 0 1 770
box -8 -3 16 105
use FILL  FILL_3741
timestamp 1711653199
transform 1 0 760 0 1 770
box -8 -3 16 105
use FILL  FILL_3742
timestamp 1711653199
transform 1 0 752 0 1 770
box -8 -3 16 105
use FILL  FILL_3743
timestamp 1711653199
transform 1 0 744 0 1 770
box -8 -3 16 105
use FILL  FILL_3744
timestamp 1711653199
transform 1 0 680 0 1 770
box -8 -3 16 105
use FILL  FILL_3745
timestamp 1711653199
transform 1 0 672 0 1 770
box -8 -3 16 105
use FILL  FILL_3746
timestamp 1711653199
transform 1 0 664 0 1 770
box -8 -3 16 105
use FILL  FILL_3747
timestamp 1711653199
transform 1 0 656 0 1 770
box -8 -3 16 105
use FILL  FILL_3748
timestamp 1711653199
transform 1 0 648 0 1 770
box -8 -3 16 105
use FILL  FILL_3749
timestamp 1711653199
transform 1 0 640 0 1 770
box -8 -3 16 105
use FILL  FILL_3750
timestamp 1711653199
transform 1 0 632 0 1 770
box -8 -3 16 105
use FILL  FILL_3751
timestamp 1711653199
transform 1 0 600 0 1 770
box -8 -3 16 105
use FILL  FILL_3752
timestamp 1711653199
transform 1 0 560 0 1 770
box -8 -3 16 105
use FILL  FILL_3753
timestamp 1711653199
transform 1 0 552 0 1 770
box -8 -3 16 105
use FILL  FILL_3754
timestamp 1711653199
transform 1 0 544 0 1 770
box -8 -3 16 105
use FILL  FILL_3755
timestamp 1711653199
transform 1 0 536 0 1 770
box -8 -3 16 105
use FILL  FILL_3756
timestamp 1711653199
transform 1 0 528 0 1 770
box -8 -3 16 105
use FILL  FILL_3757
timestamp 1711653199
transform 1 0 520 0 1 770
box -8 -3 16 105
use FILL  FILL_3758
timestamp 1711653199
transform 1 0 480 0 1 770
box -8 -3 16 105
use FILL  FILL_3759
timestamp 1711653199
transform 1 0 472 0 1 770
box -8 -3 16 105
use FILL  FILL_3760
timestamp 1711653199
transform 1 0 432 0 1 770
box -8 -3 16 105
use FILL  FILL_3761
timestamp 1711653199
transform 1 0 424 0 1 770
box -8 -3 16 105
use FILL  FILL_3762
timestamp 1711653199
transform 1 0 416 0 1 770
box -8 -3 16 105
use FILL  FILL_3763
timestamp 1711653199
transform 1 0 392 0 1 770
box -8 -3 16 105
use FILL  FILL_3764
timestamp 1711653199
transform 1 0 384 0 1 770
box -8 -3 16 105
use FILL  FILL_3765
timestamp 1711653199
transform 1 0 344 0 1 770
box -8 -3 16 105
use FILL  FILL_3766
timestamp 1711653199
transform 1 0 336 0 1 770
box -8 -3 16 105
use FILL  FILL_3767
timestamp 1711653199
transform 1 0 328 0 1 770
box -8 -3 16 105
use FILL  FILL_3768
timestamp 1711653199
transform 1 0 320 0 1 770
box -8 -3 16 105
use FILL  FILL_3769
timestamp 1711653199
transform 1 0 272 0 1 770
box -8 -3 16 105
use FILL  FILL_3770
timestamp 1711653199
transform 1 0 264 0 1 770
box -8 -3 16 105
use FILL  FILL_3771
timestamp 1711653199
transform 1 0 256 0 1 770
box -8 -3 16 105
use FILL  FILL_3772
timestamp 1711653199
transform 1 0 248 0 1 770
box -8 -3 16 105
use FILL  FILL_3773
timestamp 1711653199
transform 1 0 240 0 1 770
box -8 -3 16 105
use FILL  FILL_3774
timestamp 1711653199
transform 1 0 232 0 1 770
box -8 -3 16 105
use FILL  FILL_3775
timestamp 1711653199
transform 1 0 184 0 1 770
box -8 -3 16 105
use FILL  FILL_3776
timestamp 1711653199
transform 1 0 176 0 1 770
box -8 -3 16 105
use FILL  FILL_3777
timestamp 1711653199
transform 1 0 168 0 1 770
box -8 -3 16 105
use FILL  FILL_3778
timestamp 1711653199
transform 1 0 160 0 1 770
box -8 -3 16 105
use FILL  FILL_3779
timestamp 1711653199
transform 1 0 128 0 1 770
box -8 -3 16 105
use FILL  FILL_3780
timestamp 1711653199
transform 1 0 120 0 1 770
box -8 -3 16 105
use FILL  FILL_3781
timestamp 1711653199
transform 1 0 112 0 1 770
box -8 -3 16 105
use FILL  FILL_3782
timestamp 1711653199
transform 1 0 80 0 1 770
box -8 -3 16 105
use FILL  FILL_3783
timestamp 1711653199
transform 1 0 72 0 1 770
box -8 -3 16 105
use FILL  FILL_3784
timestamp 1711653199
transform 1 0 3392 0 -1 770
box -8 -3 16 105
use FILL  FILL_3785
timestamp 1711653199
transform 1 0 3384 0 -1 770
box -8 -3 16 105
use FILL  FILL_3786
timestamp 1711653199
transform 1 0 3376 0 -1 770
box -8 -3 16 105
use FILL  FILL_3787
timestamp 1711653199
transform 1 0 3368 0 -1 770
box -8 -3 16 105
use FILL  FILL_3788
timestamp 1711653199
transform 1 0 3360 0 -1 770
box -8 -3 16 105
use FILL  FILL_3789
timestamp 1711653199
transform 1 0 3352 0 -1 770
box -8 -3 16 105
use FILL  FILL_3790
timestamp 1711653199
transform 1 0 3344 0 -1 770
box -8 -3 16 105
use FILL  FILL_3791
timestamp 1711653199
transform 1 0 3336 0 -1 770
box -8 -3 16 105
use FILL  FILL_3792
timestamp 1711653199
transform 1 0 3328 0 -1 770
box -8 -3 16 105
use FILL  FILL_3793
timestamp 1711653199
transform 1 0 3320 0 -1 770
box -8 -3 16 105
use FILL  FILL_3794
timestamp 1711653199
transform 1 0 3272 0 -1 770
box -8 -3 16 105
use FILL  FILL_3795
timestamp 1711653199
transform 1 0 3264 0 -1 770
box -8 -3 16 105
use FILL  FILL_3796
timestamp 1711653199
transform 1 0 3256 0 -1 770
box -8 -3 16 105
use FILL  FILL_3797
timestamp 1711653199
transform 1 0 3248 0 -1 770
box -8 -3 16 105
use FILL  FILL_3798
timestamp 1711653199
transform 1 0 3240 0 -1 770
box -8 -3 16 105
use FILL  FILL_3799
timestamp 1711653199
transform 1 0 3232 0 -1 770
box -8 -3 16 105
use FILL  FILL_3800
timestamp 1711653199
transform 1 0 3224 0 -1 770
box -8 -3 16 105
use FILL  FILL_3801
timestamp 1711653199
transform 1 0 3216 0 -1 770
box -8 -3 16 105
use FILL  FILL_3802
timestamp 1711653199
transform 1 0 3208 0 -1 770
box -8 -3 16 105
use FILL  FILL_3803
timestamp 1711653199
transform 1 0 3152 0 -1 770
box -8 -3 16 105
use FILL  FILL_3804
timestamp 1711653199
transform 1 0 3144 0 -1 770
box -8 -3 16 105
use FILL  FILL_3805
timestamp 1711653199
transform 1 0 3136 0 -1 770
box -8 -3 16 105
use FILL  FILL_3806
timestamp 1711653199
transform 1 0 3128 0 -1 770
box -8 -3 16 105
use FILL  FILL_3807
timestamp 1711653199
transform 1 0 3120 0 -1 770
box -8 -3 16 105
use FILL  FILL_3808
timestamp 1711653199
transform 1 0 3112 0 -1 770
box -8 -3 16 105
use FILL  FILL_3809
timestamp 1711653199
transform 1 0 3104 0 -1 770
box -8 -3 16 105
use FILL  FILL_3810
timestamp 1711653199
transform 1 0 3064 0 -1 770
box -8 -3 16 105
use FILL  FILL_3811
timestamp 1711653199
transform 1 0 3056 0 -1 770
box -8 -3 16 105
use FILL  FILL_3812
timestamp 1711653199
transform 1 0 3032 0 -1 770
box -8 -3 16 105
use FILL  FILL_3813
timestamp 1711653199
transform 1 0 3024 0 -1 770
box -8 -3 16 105
use FILL  FILL_3814
timestamp 1711653199
transform 1 0 3016 0 -1 770
box -8 -3 16 105
use FILL  FILL_3815
timestamp 1711653199
transform 1 0 3008 0 -1 770
box -8 -3 16 105
use FILL  FILL_3816
timestamp 1711653199
transform 1 0 2968 0 -1 770
box -8 -3 16 105
use FILL  FILL_3817
timestamp 1711653199
transform 1 0 2960 0 -1 770
box -8 -3 16 105
use FILL  FILL_3818
timestamp 1711653199
transform 1 0 2952 0 -1 770
box -8 -3 16 105
use FILL  FILL_3819
timestamp 1711653199
transform 1 0 2928 0 -1 770
box -8 -3 16 105
use FILL  FILL_3820
timestamp 1711653199
transform 1 0 2920 0 -1 770
box -8 -3 16 105
use FILL  FILL_3821
timestamp 1711653199
transform 1 0 2912 0 -1 770
box -8 -3 16 105
use FILL  FILL_3822
timestamp 1711653199
transform 1 0 2904 0 -1 770
box -8 -3 16 105
use FILL  FILL_3823
timestamp 1711653199
transform 1 0 2864 0 -1 770
box -8 -3 16 105
use FILL  FILL_3824
timestamp 1711653199
transform 1 0 2856 0 -1 770
box -8 -3 16 105
use FILL  FILL_3825
timestamp 1711653199
transform 1 0 2824 0 -1 770
box -8 -3 16 105
use FILL  FILL_3826
timestamp 1711653199
transform 1 0 2816 0 -1 770
box -8 -3 16 105
use FILL  FILL_3827
timestamp 1711653199
transform 1 0 2808 0 -1 770
box -8 -3 16 105
use FILL  FILL_3828
timestamp 1711653199
transform 1 0 2800 0 -1 770
box -8 -3 16 105
use FILL  FILL_3829
timestamp 1711653199
transform 1 0 2792 0 -1 770
box -8 -3 16 105
use FILL  FILL_3830
timestamp 1711653199
transform 1 0 2728 0 -1 770
box -8 -3 16 105
use FILL  FILL_3831
timestamp 1711653199
transform 1 0 2720 0 -1 770
box -8 -3 16 105
use FILL  FILL_3832
timestamp 1711653199
transform 1 0 2712 0 -1 770
box -8 -3 16 105
use FILL  FILL_3833
timestamp 1711653199
transform 1 0 2704 0 -1 770
box -8 -3 16 105
use FILL  FILL_3834
timestamp 1711653199
transform 1 0 2696 0 -1 770
box -8 -3 16 105
use FILL  FILL_3835
timestamp 1711653199
transform 1 0 2688 0 -1 770
box -8 -3 16 105
use FILL  FILL_3836
timestamp 1711653199
transform 1 0 2648 0 -1 770
box -8 -3 16 105
use FILL  FILL_3837
timestamp 1711653199
transform 1 0 2624 0 -1 770
box -8 -3 16 105
use FILL  FILL_3838
timestamp 1711653199
transform 1 0 2616 0 -1 770
box -8 -3 16 105
use FILL  FILL_3839
timestamp 1711653199
transform 1 0 2608 0 -1 770
box -8 -3 16 105
use FILL  FILL_3840
timestamp 1711653199
transform 1 0 2600 0 -1 770
box -8 -3 16 105
use FILL  FILL_3841
timestamp 1711653199
transform 1 0 2560 0 -1 770
box -8 -3 16 105
use FILL  FILL_3842
timestamp 1711653199
transform 1 0 2552 0 -1 770
box -8 -3 16 105
use FILL  FILL_3843
timestamp 1711653199
transform 1 0 2544 0 -1 770
box -8 -3 16 105
use FILL  FILL_3844
timestamp 1711653199
transform 1 0 2536 0 -1 770
box -8 -3 16 105
use FILL  FILL_3845
timestamp 1711653199
transform 1 0 2528 0 -1 770
box -8 -3 16 105
use FILL  FILL_3846
timestamp 1711653199
transform 1 0 2520 0 -1 770
box -8 -3 16 105
use FILL  FILL_3847
timestamp 1711653199
transform 1 0 2480 0 -1 770
box -8 -3 16 105
use FILL  FILL_3848
timestamp 1711653199
transform 1 0 2472 0 -1 770
box -8 -3 16 105
use FILL  FILL_3849
timestamp 1711653199
transform 1 0 2464 0 -1 770
box -8 -3 16 105
use FILL  FILL_3850
timestamp 1711653199
transform 1 0 2456 0 -1 770
box -8 -3 16 105
use FILL  FILL_3851
timestamp 1711653199
transform 1 0 2424 0 -1 770
box -8 -3 16 105
use FILL  FILL_3852
timestamp 1711653199
transform 1 0 2416 0 -1 770
box -8 -3 16 105
use FILL  FILL_3853
timestamp 1711653199
transform 1 0 2408 0 -1 770
box -8 -3 16 105
use FILL  FILL_3854
timestamp 1711653199
transform 1 0 2400 0 -1 770
box -8 -3 16 105
use FILL  FILL_3855
timestamp 1711653199
transform 1 0 2368 0 -1 770
box -8 -3 16 105
use FILL  FILL_3856
timestamp 1711653199
transform 1 0 2360 0 -1 770
box -8 -3 16 105
use FILL  FILL_3857
timestamp 1711653199
transform 1 0 2352 0 -1 770
box -8 -3 16 105
use FILL  FILL_3858
timestamp 1711653199
transform 1 0 2320 0 -1 770
box -8 -3 16 105
use FILL  FILL_3859
timestamp 1711653199
transform 1 0 2312 0 -1 770
box -8 -3 16 105
use FILL  FILL_3860
timestamp 1711653199
transform 1 0 2304 0 -1 770
box -8 -3 16 105
use FILL  FILL_3861
timestamp 1711653199
transform 1 0 2296 0 -1 770
box -8 -3 16 105
use FILL  FILL_3862
timestamp 1711653199
transform 1 0 2288 0 -1 770
box -8 -3 16 105
use FILL  FILL_3863
timestamp 1711653199
transform 1 0 2256 0 -1 770
box -8 -3 16 105
use FILL  FILL_3864
timestamp 1711653199
transform 1 0 2248 0 -1 770
box -8 -3 16 105
use FILL  FILL_3865
timestamp 1711653199
transform 1 0 2208 0 -1 770
box -8 -3 16 105
use FILL  FILL_3866
timestamp 1711653199
transform 1 0 2200 0 -1 770
box -8 -3 16 105
use FILL  FILL_3867
timestamp 1711653199
transform 1 0 2192 0 -1 770
box -8 -3 16 105
use FILL  FILL_3868
timestamp 1711653199
transform 1 0 2184 0 -1 770
box -8 -3 16 105
use FILL  FILL_3869
timestamp 1711653199
transform 1 0 2144 0 -1 770
box -8 -3 16 105
use FILL  FILL_3870
timestamp 1711653199
transform 1 0 2136 0 -1 770
box -8 -3 16 105
use FILL  FILL_3871
timestamp 1711653199
transform 1 0 2128 0 -1 770
box -8 -3 16 105
use FILL  FILL_3872
timestamp 1711653199
transform 1 0 2120 0 -1 770
box -8 -3 16 105
use FILL  FILL_3873
timestamp 1711653199
transform 1 0 2088 0 -1 770
box -8 -3 16 105
use FILL  FILL_3874
timestamp 1711653199
transform 1 0 2080 0 -1 770
box -8 -3 16 105
use FILL  FILL_3875
timestamp 1711653199
transform 1 0 2072 0 -1 770
box -8 -3 16 105
use FILL  FILL_3876
timestamp 1711653199
transform 1 0 2064 0 -1 770
box -8 -3 16 105
use FILL  FILL_3877
timestamp 1711653199
transform 1 0 2056 0 -1 770
box -8 -3 16 105
use FILL  FILL_3878
timestamp 1711653199
transform 1 0 2048 0 -1 770
box -8 -3 16 105
use FILL  FILL_3879
timestamp 1711653199
transform 1 0 2000 0 -1 770
box -8 -3 16 105
use FILL  FILL_3880
timestamp 1711653199
transform 1 0 1992 0 -1 770
box -8 -3 16 105
use FILL  FILL_3881
timestamp 1711653199
transform 1 0 1984 0 -1 770
box -8 -3 16 105
use FILL  FILL_3882
timestamp 1711653199
transform 1 0 1976 0 -1 770
box -8 -3 16 105
use FILL  FILL_3883
timestamp 1711653199
transform 1 0 1968 0 -1 770
box -8 -3 16 105
use FILL  FILL_3884
timestamp 1711653199
transform 1 0 1936 0 -1 770
box -8 -3 16 105
use FILL  FILL_3885
timestamp 1711653199
transform 1 0 1928 0 -1 770
box -8 -3 16 105
use FILL  FILL_3886
timestamp 1711653199
transform 1 0 1920 0 -1 770
box -8 -3 16 105
use FILL  FILL_3887
timestamp 1711653199
transform 1 0 1912 0 -1 770
box -8 -3 16 105
use FILL  FILL_3888
timestamp 1711653199
transform 1 0 1904 0 -1 770
box -8 -3 16 105
use FILL  FILL_3889
timestamp 1711653199
transform 1 0 1896 0 -1 770
box -8 -3 16 105
use FILL  FILL_3890
timestamp 1711653199
transform 1 0 1848 0 -1 770
box -8 -3 16 105
use FILL  FILL_3891
timestamp 1711653199
transform 1 0 1840 0 -1 770
box -8 -3 16 105
use FILL  FILL_3892
timestamp 1711653199
transform 1 0 1832 0 -1 770
box -8 -3 16 105
use FILL  FILL_3893
timestamp 1711653199
transform 1 0 1824 0 -1 770
box -8 -3 16 105
use FILL  FILL_3894
timestamp 1711653199
transform 1 0 1816 0 -1 770
box -8 -3 16 105
use FILL  FILL_3895
timestamp 1711653199
transform 1 0 1784 0 -1 770
box -8 -3 16 105
use FILL  FILL_3896
timestamp 1711653199
transform 1 0 1776 0 -1 770
box -8 -3 16 105
use FILL  FILL_3897
timestamp 1711653199
transform 1 0 1768 0 -1 770
box -8 -3 16 105
use FILL  FILL_3898
timestamp 1711653199
transform 1 0 1744 0 -1 770
box -8 -3 16 105
use FILL  FILL_3899
timestamp 1711653199
transform 1 0 1736 0 -1 770
box -8 -3 16 105
use FILL  FILL_3900
timestamp 1711653199
transform 1 0 1728 0 -1 770
box -8 -3 16 105
use FILL  FILL_3901
timestamp 1711653199
transform 1 0 1720 0 -1 770
box -8 -3 16 105
use FILL  FILL_3902
timestamp 1711653199
transform 1 0 1696 0 -1 770
box -8 -3 16 105
use FILL  FILL_3903
timestamp 1711653199
transform 1 0 1688 0 -1 770
box -8 -3 16 105
use FILL  FILL_3904
timestamp 1711653199
transform 1 0 1680 0 -1 770
box -8 -3 16 105
use FILL  FILL_3905
timestamp 1711653199
transform 1 0 1672 0 -1 770
box -8 -3 16 105
use FILL  FILL_3906
timestamp 1711653199
transform 1 0 1632 0 -1 770
box -8 -3 16 105
use FILL  FILL_3907
timestamp 1711653199
transform 1 0 1624 0 -1 770
box -8 -3 16 105
use FILL  FILL_3908
timestamp 1711653199
transform 1 0 1616 0 -1 770
box -8 -3 16 105
use FILL  FILL_3909
timestamp 1711653199
transform 1 0 1608 0 -1 770
box -8 -3 16 105
use FILL  FILL_3910
timestamp 1711653199
transform 1 0 1600 0 -1 770
box -8 -3 16 105
use FILL  FILL_3911
timestamp 1711653199
transform 1 0 1592 0 -1 770
box -8 -3 16 105
use FILL  FILL_3912
timestamp 1711653199
transform 1 0 1584 0 -1 770
box -8 -3 16 105
use FILL  FILL_3913
timestamp 1711653199
transform 1 0 1552 0 -1 770
box -8 -3 16 105
use FILL  FILL_3914
timestamp 1711653199
transform 1 0 1544 0 -1 770
box -8 -3 16 105
use FILL  FILL_3915
timestamp 1711653199
transform 1 0 1512 0 -1 770
box -8 -3 16 105
use FILL  FILL_3916
timestamp 1711653199
transform 1 0 1504 0 -1 770
box -8 -3 16 105
use FILL  FILL_3917
timestamp 1711653199
transform 1 0 1496 0 -1 770
box -8 -3 16 105
use FILL  FILL_3918
timestamp 1711653199
transform 1 0 1488 0 -1 770
box -8 -3 16 105
use FILL  FILL_3919
timestamp 1711653199
transform 1 0 1480 0 -1 770
box -8 -3 16 105
use FILL  FILL_3920
timestamp 1711653199
transform 1 0 1472 0 -1 770
box -8 -3 16 105
use FILL  FILL_3921
timestamp 1711653199
transform 1 0 1424 0 -1 770
box -8 -3 16 105
use FILL  FILL_3922
timestamp 1711653199
transform 1 0 1416 0 -1 770
box -8 -3 16 105
use FILL  FILL_3923
timestamp 1711653199
transform 1 0 1408 0 -1 770
box -8 -3 16 105
use FILL  FILL_3924
timestamp 1711653199
transform 1 0 1400 0 -1 770
box -8 -3 16 105
use FILL  FILL_3925
timestamp 1711653199
transform 1 0 1392 0 -1 770
box -8 -3 16 105
use FILL  FILL_3926
timestamp 1711653199
transform 1 0 1384 0 -1 770
box -8 -3 16 105
use FILL  FILL_3927
timestamp 1711653199
transform 1 0 1352 0 -1 770
box -8 -3 16 105
use FILL  FILL_3928
timestamp 1711653199
transform 1 0 1344 0 -1 770
box -8 -3 16 105
use FILL  FILL_3929
timestamp 1711653199
transform 1 0 1336 0 -1 770
box -8 -3 16 105
use FILL  FILL_3930
timestamp 1711653199
transform 1 0 1304 0 -1 770
box -8 -3 16 105
use FILL  FILL_3931
timestamp 1711653199
transform 1 0 1296 0 -1 770
box -8 -3 16 105
use FILL  FILL_3932
timestamp 1711653199
transform 1 0 1288 0 -1 770
box -8 -3 16 105
use FILL  FILL_3933
timestamp 1711653199
transform 1 0 1280 0 -1 770
box -8 -3 16 105
use FILL  FILL_3934
timestamp 1711653199
transform 1 0 1272 0 -1 770
box -8 -3 16 105
use FILL  FILL_3935
timestamp 1711653199
transform 1 0 1248 0 -1 770
box -8 -3 16 105
use FILL  FILL_3936
timestamp 1711653199
transform 1 0 1240 0 -1 770
box -8 -3 16 105
use FILL  FILL_3937
timestamp 1711653199
transform 1 0 1232 0 -1 770
box -8 -3 16 105
use FILL  FILL_3938
timestamp 1711653199
transform 1 0 1200 0 -1 770
box -8 -3 16 105
use FILL  FILL_3939
timestamp 1711653199
transform 1 0 1192 0 -1 770
box -8 -3 16 105
use FILL  FILL_3940
timestamp 1711653199
transform 1 0 1184 0 -1 770
box -8 -3 16 105
use FILL  FILL_3941
timestamp 1711653199
transform 1 0 1176 0 -1 770
box -8 -3 16 105
use FILL  FILL_3942
timestamp 1711653199
transform 1 0 1168 0 -1 770
box -8 -3 16 105
use FILL  FILL_3943
timestamp 1711653199
transform 1 0 1160 0 -1 770
box -8 -3 16 105
use FILL  FILL_3944
timestamp 1711653199
transform 1 0 1112 0 -1 770
box -8 -3 16 105
use FILL  FILL_3945
timestamp 1711653199
transform 1 0 1104 0 -1 770
box -8 -3 16 105
use FILL  FILL_3946
timestamp 1711653199
transform 1 0 1096 0 -1 770
box -8 -3 16 105
use FILL  FILL_3947
timestamp 1711653199
transform 1 0 1088 0 -1 770
box -8 -3 16 105
use FILL  FILL_3948
timestamp 1711653199
transform 1 0 1048 0 -1 770
box -8 -3 16 105
use FILL  FILL_3949
timestamp 1711653199
transform 1 0 1040 0 -1 770
box -8 -3 16 105
use FILL  FILL_3950
timestamp 1711653199
transform 1 0 1032 0 -1 770
box -8 -3 16 105
use FILL  FILL_3951
timestamp 1711653199
transform 1 0 1000 0 -1 770
box -8 -3 16 105
use FILL  FILL_3952
timestamp 1711653199
transform 1 0 992 0 -1 770
box -8 -3 16 105
use FILL  FILL_3953
timestamp 1711653199
transform 1 0 968 0 -1 770
box -8 -3 16 105
use FILL  FILL_3954
timestamp 1711653199
transform 1 0 944 0 -1 770
box -8 -3 16 105
use FILL  FILL_3955
timestamp 1711653199
transform 1 0 936 0 -1 770
box -8 -3 16 105
use FILL  FILL_3956
timestamp 1711653199
transform 1 0 928 0 -1 770
box -8 -3 16 105
use FILL  FILL_3957
timestamp 1711653199
transform 1 0 920 0 -1 770
box -8 -3 16 105
use FILL  FILL_3958
timestamp 1711653199
transform 1 0 872 0 -1 770
box -8 -3 16 105
use FILL  FILL_3959
timestamp 1711653199
transform 1 0 864 0 -1 770
box -8 -3 16 105
use FILL  FILL_3960
timestamp 1711653199
transform 1 0 856 0 -1 770
box -8 -3 16 105
use FILL  FILL_3961
timestamp 1711653199
transform 1 0 848 0 -1 770
box -8 -3 16 105
use FILL  FILL_3962
timestamp 1711653199
transform 1 0 808 0 -1 770
box -8 -3 16 105
use FILL  FILL_3963
timestamp 1711653199
transform 1 0 800 0 -1 770
box -8 -3 16 105
use FILL  FILL_3964
timestamp 1711653199
transform 1 0 792 0 -1 770
box -8 -3 16 105
use FILL  FILL_3965
timestamp 1711653199
transform 1 0 744 0 -1 770
box -8 -3 16 105
use FILL  FILL_3966
timestamp 1711653199
transform 1 0 736 0 -1 770
box -8 -3 16 105
use FILL  FILL_3967
timestamp 1711653199
transform 1 0 728 0 -1 770
box -8 -3 16 105
use FILL  FILL_3968
timestamp 1711653199
transform 1 0 720 0 -1 770
box -8 -3 16 105
use FILL  FILL_3969
timestamp 1711653199
transform 1 0 712 0 -1 770
box -8 -3 16 105
use FILL  FILL_3970
timestamp 1711653199
transform 1 0 656 0 -1 770
box -8 -3 16 105
use FILL  FILL_3971
timestamp 1711653199
transform 1 0 648 0 -1 770
box -8 -3 16 105
use FILL  FILL_3972
timestamp 1711653199
transform 1 0 640 0 -1 770
box -8 -3 16 105
use FILL  FILL_3973
timestamp 1711653199
transform 1 0 632 0 -1 770
box -8 -3 16 105
use FILL  FILL_3974
timestamp 1711653199
transform 1 0 560 0 -1 770
box -8 -3 16 105
use FILL  FILL_3975
timestamp 1711653199
transform 1 0 552 0 -1 770
box -8 -3 16 105
use FILL  FILL_3976
timestamp 1711653199
transform 1 0 544 0 -1 770
box -8 -3 16 105
use FILL  FILL_3977
timestamp 1711653199
transform 1 0 536 0 -1 770
box -8 -3 16 105
use FILL  FILL_3978
timestamp 1711653199
transform 1 0 528 0 -1 770
box -8 -3 16 105
use FILL  FILL_3979
timestamp 1711653199
transform 1 0 464 0 -1 770
box -8 -3 16 105
use FILL  FILL_3980
timestamp 1711653199
transform 1 0 456 0 -1 770
box -8 -3 16 105
use FILL  FILL_3981
timestamp 1711653199
transform 1 0 448 0 -1 770
box -8 -3 16 105
use FILL  FILL_3982
timestamp 1711653199
transform 1 0 440 0 -1 770
box -8 -3 16 105
use FILL  FILL_3983
timestamp 1711653199
transform 1 0 432 0 -1 770
box -8 -3 16 105
use FILL  FILL_3984
timestamp 1711653199
transform 1 0 384 0 -1 770
box -8 -3 16 105
use FILL  FILL_3985
timestamp 1711653199
transform 1 0 352 0 -1 770
box -8 -3 16 105
use FILL  FILL_3986
timestamp 1711653199
transform 1 0 344 0 -1 770
box -8 -3 16 105
use FILL  FILL_3987
timestamp 1711653199
transform 1 0 336 0 -1 770
box -8 -3 16 105
use FILL  FILL_3988
timestamp 1711653199
transform 1 0 328 0 -1 770
box -8 -3 16 105
use FILL  FILL_3989
timestamp 1711653199
transform 1 0 288 0 -1 770
box -8 -3 16 105
use FILL  FILL_3990
timestamp 1711653199
transform 1 0 280 0 -1 770
box -8 -3 16 105
use FILL  FILL_3991
timestamp 1711653199
transform 1 0 272 0 -1 770
box -8 -3 16 105
use FILL  FILL_3992
timestamp 1711653199
transform 1 0 264 0 -1 770
box -8 -3 16 105
use FILL  FILL_3993
timestamp 1711653199
transform 1 0 216 0 -1 770
box -8 -3 16 105
use FILL  FILL_3994
timestamp 1711653199
transform 1 0 208 0 -1 770
box -8 -3 16 105
use FILL  FILL_3995
timestamp 1711653199
transform 1 0 200 0 -1 770
box -8 -3 16 105
use FILL  FILL_3996
timestamp 1711653199
transform 1 0 192 0 -1 770
box -8 -3 16 105
use FILL  FILL_3997
timestamp 1711653199
transform 1 0 152 0 -1 770
box -8 -3 16 105
use FILL  FILL_3998
timestamp 1711653199
transform 1 0 144 0 -1 770
box -8 -3 16 105
use FILL  FILL_3999
timestamp 1711653199
transform 1 0 136 0 -1 770
box -8 -3 16 105
use FILL  FILL_4000
timestamp 1711653199
transform 1 0 128 0 -1 770
box -8 -3 16 105
use FILL  FILL_4001
timestamp 1711653199
transform 1 0 80 0 -1 770
box -8 -3 16 105
use FILL  FILL_4002
timestamp 1711653199
transform 1 0 72 0 -1 770
box -8 -3 16 105
use FILL  FILL_4003
timestamp 1711653199
transform 1 0 3392 0 1 570
box -8 -3 16 105
use FILL  FILL_4004
timestamp 1711653199
transform 1 0 3384 0 1 570
box -8 -3 16 105
use FILL  FILL_4005
timestamp 1711653199
transform 1 0 3360 0 1 570
box -8 -3 16 105
use FILL  FILL_4006
timestamp 1711653199
transform 1 0 3320 0 1 570
box -8 -3 16 105
use FILL  FILL_4007
timestamp 1711653199
transform 1 0 3312 0 1 570
box -8 -3 16 105
use FILL  FILL_4008
timestamp 1711653199
transform 1 0 3272 0 1 570
box -8 -3 16 105
use FILL  FILL_4009
timestamp 1711653199
transform 1 0 3264 0 1 570
box -8 -3 16 105
use FILL  FILL_4010
timestamp 1711653199
transform 1 0 3256 0 1 570
box -8 -3 16 105
use FILL  FILL_4011
timestamp 1711653199
transform 1 0 3224 0 1 570
box -8 -3 16 105
use FILL  FILL_4012
timestamp 1711653199
transform 1 0 3216 0 1 570
box -8 -3 16 105
use FILL  FILL_4013
timestamp 1711653199
transform 1 0 3208 0 1 570
box -8 -3 16 105
use FILL  FILL_4014
timestamp 1711653199
transform 1 0 3200 0 1 570
box -8 -3 16 105
use FILL  FILL_4015
timestamp 1711653199
transform 1 0 3192 0 1 570
box -8 -3 16 105
use FILL  FILL_4016
timestamp 1711653199
transform 1 0 3160 0 1 570
box -8 -3 16 105
use FILL  FILL_4017
timestamp 1711653199
transform 1 0 3152 0 1 570
box -8 -3 16 105
use FILL  FILL_4018
timestamp 1711653199
transform 1 0 3144 0 1 570
box -8 -3 16 105
use FILL  FILL_4019
timestamp 1711653199
transform 1 0 3136 0 1 570
box -8 -3 16 105
use FILL  FILL_4020
timestamp 1711653199
transform 1 0 3104 0 1 570
box -8 -3 16 105
use FILL  FILL_4021
timestamp 1711653199
transform 1 0 3096 0 1 570
box -8 -3 16 105
use FILL  FILL_4022
timestamp 1711653199
transform 1 0 3088 0 1 570
box -8 -3 16 105
use FILL  FILL_4023
timestamp 1711653199
transform 1 0 3080 0 1 570
box -8 -3 16 105
use FILL  FILL_4024
timestamp 1711653199
transform 1 0 3072 0 1 570
box -8 -3 16 105
use FILL  FILL_4025
timestamp 1711653199
transform 1 0 3032 0 1 570
box -8 -3 16 105
use FILL  FILL_4026
timestamp 1711653199
transform 1 0 3024 0 1 570
box -8 -3 16 105
use FILL  FILL_4027
timestamp 1711653199
transform 1 0 3016 0 1 570
box -8 -3 16 105
use FILL  FILL_4028
timestamp 1711653199
transform 1 0 3008 0 1 570
box -8 -3 16 105
use FILL  FILL_4029
timestamp 1711653199
transform 1 0 3000 0 1 570
box -8 -3 16 105
use FILL  FILL_4030
timestamp 1711653199
transform 1 0 2992 0 1 570
box -8 -3 16 105
use FILL  FILL_4031
timestamp 1711653199
transform 1 0 2984 0 1 570
box -8 -3 16 105
use FILL  FILL_4032
timestamp 1711653199
transform 1 0 2928 0 1 570
box -8 -3 16 105
use FILL  FILL_4033
timestamp 1711653199
transform 1 0 2920 0 1 570
box -8 -3 16 105
use FILL  FILL_4034
timestamp 1711653199
transform 1 0 2912 0 1 570
box -8 -3 16 105
use FILL  FILL_4035
timestamp 1711653199
transform 1 0 2904 0 1 570
box -8 -3 16 105
use FILL  FILL_4036
timestamp 1711653199
transform 1 0 2896 0 1 570
box -8 -3 16 105
use FILL  FILL_4037
timestamp 1711653199
transform 1 0 2888 0 1 570
box -8 -3 16 105
use FILL  FILL_4038
timestamp 1711653199
transform 1 0 2880 0 1 570
box -8 -3 16 105
use FILL  FILL_4039
timestamp 1711653199
transform 1 0 2832 0 1 570
box -8 -3 16 105
use FILL  FILL_4040
timestamp 1711653199
transform 1 0 2824 0 1 570
box -8 -3 16 105
use FILL  FILL_4041
timestamp 1711653199
transform 1 0 2816 0 1 570
box -8 -3 16 105
use FILL  FILL_4042
timestamp 1711653199
transform 1 0 2776 0 1 570
box -8 -3 16 105
use FILL  FILL_4043
timestamp 1711653199
transform 1 0 2768 0 1 570
box -8 -3 16 105
use FILL  FILL_4044
timestamp 1711653199
transform 1 0 2760 0 1 570
box -8 -3 16 105
use FILL  FILL_4045
timestamp 1711653199
transform 1 0 2728 0 1 570
box -8 -3 16 105
use FILL  FILL_4046
timestamp 1711653199
transform 1 0 2720 0 1 570
box -8 -3 16 105
use FILL  FILL_4047
timestamp 1711653199
transform 1 0 2712 0 1 570
box -8 -3 16 105
use FILL  FILL_4048
timestamp 1711653199
transform 1 0 2664 0 1 570
box -8 -3 16 105
use FILL  FILL_4049
timestamp 1711653199
transform 1 0 2656 0 1 570
box -8 -3 16 105
use FILL  FILL_4050
timestamp 1711653199
transform 1 0 2648 0 1 570
box -8 -3 16 105
use FILL  FILL_4051
timestamp 1711653199
transform 1 0 2640 0 1 570
box -8 -3 16 105
use FILL  FILL_4052
timestamp 1711653199
transform 1 0 2632 0 1 570
box -8 -3 16 105
use FILL  FILL_4053
timestamp 1711653199
transform 1 0 2592 0 1 570
box -8 -3 16 105
use FILL  FILL_4054
timestamp 1711653199
transform 1 0 2584 0 1 570
box -8 -3 16 105
use FILL  FILL_4055
timestamp 1711653199
transform 1 0 2576 0 1 570
box -8 -3 16 105
use FILL  FILL_4056
timestamp 1711653199
transform 1 0 2568 0 1 570
box -8 -3 16 105
use FILL  FILL_4057
timestamp 1711653199
transform 1 0 2520 0 1 570
box -8 -3 16 105
use FILL  FILL_4058
timestamp 1711653199
transform 1 0 2512 0 1 570
box -8 -3 16 105
use FILL  FILL_4059
timestamp 1711653199
transform 1 0 2504 0 1 570
box -8 -3 16 105
use FILL  FILL_4060
timestamp 1711653199
transform 1 0 2496 0 1 570
box -8 -3 16 105
use FILL  FILL_4061
timestamp 1711653199
transform 1 0 2488 0 1 570
box -8 -3 16 105
use FILL  FILL_4062
timestamp 1711653199
transform 1 0 2448 0 1 570
box -8 -3 16 105
use FILL  FILL_4063
timestamp 1711653199
transform 1 0 2440 0 1 570
box -8 -3 16 105
use FILL  FILL_4064
timestamp 1711653199
transform 1 0 2432 0 1 570
box -8 -3 16 105
use FILL  FILL_4065
timestamp 1711653199
transform 1 0 2424 0 1 570
box -8 -3 16 105
use FILL  FILL_4066
timestamp 1711653199
transform 1 0 2416 0 1 570
box -8 -3 16 105
use FILL  FILL_4067
timestamp 1711653199
transform 1 0 2376 0 1 570
box -8 -3 16 105
use FILL  FILL_4068
timestamp 1711653199
transform 1 0 2344 0 1 570
box -8 -3 16 105
use FILL  FILL_4069
timestamp 1711653199
transform 1 0 2336 0 1 570
box -8 -3 16 105
use FILL  FILL_4070
timestamp 1711653199
transform 1 0 2328 0 1 570
box -8 -3 16 105
use FILL  FILL_4071
timestamp 1711653199
transform 1 0 2320 0 1 570
box -8 -3 16 105
use FILL  FILL_4072
timestamp 1711653199
transform 1 0 2312 0 1 570
box -8 -3 16 105
use FILL  FILL_4073
timestamp 1711653199
transform 1 0 2304 0 1 570
box -8 -3 16 105
use FILL  FILL_4074
timestamp 1711653199
transform 1 0 2296 0 1 570
box -8 -3 16 105
use FILL  FILL_4075
timestamp 1711653199
transform 1 0 2248 0 1 570
box -8 -3 16 105
use FILL  FILL_4076
timestamp 1711653199
transform 1 0 2240 0 1 570
box -8 -3 16 105
use FILL  FILL_4077
timestamp 1711653199
transform 1 0 2232 0 1 570
box -8 -3 16 105
use FILL  FILL_4078
timestamp 1711653199
transform 1 0 2224 0 1 570
box -8 -3 16 105
use FILL  FILL_4079
timestamp 1711653199
transform 1 0 2184 0 1 570
box -8 -3 16 105
use FILL  FILL_4080
timestamp 1711653199
transform 1 0 2176 0 1 570
box -8 -3 16 105
use FILL  FILL_4081
timestamp 1711653199
transform 1 0 2168 0 1 570
box -8 -3 16 105
use FILL  FILL_4082
timestamp 1711653199
transform 1 0 2128 0 1 570
box -8 -3 16 105
use FILL  FILL_4083
timestamp 1711653199
transform 1 0 2120 0 1 570
box -8 -3 16 105
use FILL  FILL_4084
timestamp 1711653199
transform 1 0 2112 0 1 570
box -8 -3 16 105
use FILL  FILL_4085
timestamp 1711653199
transform 1 0 2104 0 1 570
box -8 -3 16 105
use FILL  FILL_4086
timestamp 1711653199
transform 1 0 2064 0 1 570
box -8 -3 16 105
use FILL  FILL_4087
timestamp 1711653199
transform 1 0 2056 0 1 570
box -8 -3 16 105
use FILL  FILL_4088
timestamp 1711653199
transform 1 0 2048 0 1 570
box -8 -3 16 105
use FILL  FILL_4089
timestamp 1711653199
transform 1 0 2040 0 1 570
box -8 -3 16 105
use FILL  FILL_4090
timestamp 1711653199
transform 1 0 2000 0 1 570
box -8 -3 16 105
use FILL  FILL_4091
timestamp 1711653199
transform 1 0 1992 0 1 570
box -8 -3 16 105
use FILL  FILL_4092
timestamp 1711653199
transform 1 0 1984 0 1 570
box -8 -3 16 105
use FILL  FILL_4093
timestamp 1711653199
transform 1 0 1976 0 1 570
box -8 -3 16 105
use FILL  FILL_4094
timestamp 1711653199
transform 1 0 1968 0 1 570
box -8 -3 16 105
use FILL  FILL_4095
timestamp 1711653199
transform 1 0 1960 0 1 570
box -8 -3 16 105
use FILL  FILL_4096
timestamp 1711653199
transform 1 0 1912 0 1 570
box -8 -3 16 105
use FILL  FILL_4097
timestamp 1711653199
transform 1 0 1904 0 1 570
box -8 -3 16 105
use FILL  FILL_4098
timestamp 1711653199
transform 1 0 1896 0 1 570
box -8 -3 16 105
use FILL  FILL_4099
timestamp 1711653199
transform 1 0 1888 0 1 570
box -8 -3 16 105
use FILL  FILL_4100
timestamp 1711653199
transform 1 0 1880 0 1 570
box -8 -3 16 105
use FILL  FILL_4101
timestamp 1711653199
transform 1 0 1872 0 1 570
box -8 -3 16 105
use FILL  FILL_4102
timestamp 1711653199
transform 1 0 1832 0 1 570
box -8 -3 16 105
use FILL  FILL_4103
timestamp 1711653199
transform 1 0 1824 0 1 570
box -8 -3 16 105
use FILL  FILL_4104
timestamp 1711653199
transform 1 0 1816 0 1 570
box -8 -3 16 105
use FILL  FILL_4105
timestamp 1711653199
transform 1 0 1784 0 1 570
box -8 -3 16 105
use FILL  FILL_4106
timestamp 1711653199
transform 1 0 1776 0 1 570
box -8 -3 16 105
use FILL  FILL_4107
timestamp 1711653199
transform 1 0 1768 0 1 570
box -8 -3 16 105
use FILL  FILL_4108
timestamp 1711653199
transform 1 0 1760 0 1 570
box -8 -3 16 105
use FILL  FILL_4109
timestamp 1711653199
transform 1 0 1752 0 1 570
box -8 -3 16 105
use FILL  FILL_4110
timestamp 1711653199
transform 1 0 1744 0 1 570
box -8 -3 16 105
use FILL  FILL_4111
timestamp 1711653199
transform 1 0 1704 0 1 570
box -8 -3 16 105
use FILL  FILL_4112
timestamp 1711653199
transform 1 0 1696 0 1 570
box -8 -3 16 105
use FILL  FILL_4113
timestamp 1711653199
transform 1 0 1688 0 1 570
box -8 -3 16 105
use FILL  FILL_4114
timestamp 1711653199
transform 1 0 1680 0 1 570
box -8 -3 16 105
use FILL  FILL_4115
timestamp 1711653199
transform 1 0 1672 0 1 570
box -8 -3 16 105
use FILL  FILL_4116
timestamp 1711653199
transform 1 0 1648 0 1 570
box -8 -3 16 105
use FILL  FILL_4117
timestamp 1711653199
transform 1 0 1640 0 1 570
box -8 -3 16 105
use FILL  FILL_4118
timestamp 1711653199
transform 1 0 1632 0 1 570
box -8 -3 16 105
use FILL  FILL_4119
timestamp 1711653199
transform 1 0 1624 0 1 570
box -8 -3 16 105
use FILL  FILL_4120
timestamp 1711653199
transform 1 0 1584 0 1 570
box -8 -3 16 105
use FILL  FILL_4121
timestamp 1711653199
transform 1 0 1576 0 1 570
box -8 -3 16 105
use FILL  FILL_4122
timestamp 1711653199
transform 1 0 1568 0 1 570
box -8 -3 16 105
use FILL  FILL_4123
timestamp 1711653199
transform 1 0 1560 0 1 570
box -8 -3 16 105
use FILL  FILL_4124
timestamp 1711653199
transform 1 0 1552 0 1 570
box -8 -3 16 105
use FILL  FILL_4125
timestamp 1711653199
transform 1 0 1544 0 1 570
box -8 -3 16 105
use FILL  FILL_4126
timestamp 1711653199
transform 1 0 1536 0 1 570
box -8 -3 16 105
use FILL  FILL_4127
timestamp 1711653199
transform 1 0 1488 0 1 570
box -8 -3 16 105
use FILL  FILL_4128
timestamp 1711653199
transform 1 0 1480 0 1 570
box -8 -3 16 105
use FILL  FILL_4129
timestamp 1711653199
transform 1 0 1472 0 1 570
box -8 -3 16 105
use FILL  FILL_4130
timestamp 1711653199
transform 1 0 1464 0 1 570
box -8 -3 16 105
use FILL  FILL_4131
timestamp 1711653199
transform 1 0 1456 0 1 570
box -8 -3 16 105
use FILL  FILL_4132
timestamp 1711653199
transform 1 0 1448 0 1 570
box -8 -3 16 105
use FILL  FILL_4133
timestamp 1711653199
transform 1 0 1408 0 1 570
box -8 -3 16 105
use FILL  FILL_4134
timestamp 1711653199
transform 1 0 1400 0 1 570
box -8 -3 16 105
use FILL  FILL_4135
timestamp 1711653199
transform 1 0 1392 0 1 570
box -8 -3 16 105
use FILL  FILL_4136
timestamp 1711653199
transform 1 0 1384 0 1 570
box -8 -3 16 105
use FILL  FILL_4137
timestamp 1711653199
transform 1 0 1376 0 1 570
box -8 -3 16 105
use FILL  FILL_4138
timestamp 1711653199
transform 1 0 1336 0 1 570
box -8 -3 16 105
use FILL  FILL_4139
timestamp 1711653199
transform 1 0 1328 0 1 570
box -8 -3 16 105
use FILL  FILL_4140
timestamp 1711653199
transform 1 0 1320 0 1 570
box -8 -3 16 105
use FILL  FILL_4141
timestamp 1711653199
transform 1 0 1312 0 1 570
box -8 -3 16 105
use FILL  FILL_4142
timestamp 1711653199
transform 1 0 1264 0 1 570
box -8 -3 16 105
use FILL  FILL_4143
timestamp 1711653199
transform 1 0 1256 0 1 570
box -8 -3 16 105
use FILL  FILL_4144
timestamp 1711653199
transform 1 0 1248 0 1 570
box -8 -3 16 105
use FILL  FILL_4145
timestamp 1711653199
transform 1 0 1240 0 1 570
box -8 -3 16 105
use FILL  FILL_4146
timestamp 1711653199
transform 1 0 1232 0 1 570
box -8 -3 16 105
use FILL  FILL_4147
timestamp 1711653199
transform 1 0 1224 0 1 570
box -8 -3 16 105
use FILL  FILL_4148
timestamp 1711653199
transform 1 0 1184 0 1 570
box -8 -3 16 105
use FILL  FILL_4149
timestamp 1711653199
transform 1 0 1176 0 1 570
box -8 -3 16 105
use FILL  FILL_4150
timestamp 1711653199
transform 1 0 1168 0 1 570
box -8 -3 16 105
use FILL  FILL_4151
timestamp 1711653199
transform 1 0 1128 0 1 570
box -8 -3 16 105
use FILL  FILL_4152
timestamp 1711653199
transform 1 0 1120 0 1 570
box -8 -3 16 105
use FILL  FILL_4153
timestamp 1711653199
transform 1 0 1112 0 1 570
box -8 -3 16 105
use FILL  FILL_4154
timestamp 1711653199
transform 1 0 1072 0 1 570
box -8 -3 16 105
use FILL  FILL_4155
timestamp 1711653199
transform 1 0 1064 0 1 570
box -8 -3 16 105
use FILL  FILL_4156
timestamp 1711653199
transform 1 0 1056 0 1 570
box -8 -3 16 105
use FILL  FILL_4157
timestamp 1711653199
transform 1 0 1016 0 1 570
box -8 -3 16 105
use FILL  FILL_4158
timestamp 1711653199
transform 1 0 1008 0 1 570
box -8 -3 16 105
use FILL  FILL_4159
timestamp 1711653199
transform 1 0 1000 0 1 570
box -8 -3 16 105
use FILL  FILL_4160
timestamp 1711653199
transform 1 0 992 0 1 570
box -8 -3 16 105
use FILL  FILL_4161
timestamp 1711653199
transform 1 0 984 0 1 570
box -8 -3 16 105
use FILL  FILL_4162
timestamp 1711653199
transform 1 0 976 0 1 570
box -8 -3 16 105
use FILL  FILL_4163
timestamp 1711653199
transform 1 0 928 0 1 570
box -8 -3 16 105
use FILL  FILL_4164
timestamp 1711653199
transform 1 0 920 0 1 570
box -8 -3 16 105
use FILL  FILL_4165
timestamp 1711653199
transform 1 0 912 0 1 570
box -8 -3 16 105
use FILL  FILL_4166
timestamp 1711653199
transform 1 0 904 0 1 570
box -8 -3 16 105
use FILL  FILL_4167
timestamp 1711653199
transform 1 0 896 0 1 570
box -8 -3 16 105
use FILL  FILL_4168
timestamp 1711653199
transform 1 0 864 0 1 570
box -8 -3 16 105
use FILL  FILL_4169
timestamp 1711653199
transform 1 0 856 0 1 570
box -8 -3 16 105
use FILL  FILL_4170
timestamp 1711653199
transform 1 0 848 0 1 570
box -8 -3 16 105
use FILL  FILL_4171
timestamp 1711653199
transform 1 0 808 0 1 570
box -8 -3 16 105
use FILL  FILL_4172
timestamp 1711653199
transform 1 0 800 0 1 570
box -8 -3 16 105
use FILL  FILL_4173
timestamp 1711653199
transform 1 0 792 0 1 570
box -8 -3 16 105
use FILL  FILL_4174
timestamp 1711653199
transform 1 0 784 0 1 570
box -8 -3 16 105
use FILL  FILL_4175
timestamp 1711653199
transform 1 0 752 0 1 570
box -8 -3 16 105
use FILL  FILL_4176
timestamp 1711653199
transform 1 0 744 0 1 570
box -8 -3 16 105
use FILL  FILL_4177
timestamp 1711653199
transform 1 0 736 0 1 570
box -8 -3 16 105
use FILL  FILL_4178
timestamp 1711653199
transform 1 0 704 0 1 570
box -8 -3 16 105
use FILL  FILL_4179
timestamp 1711653199
transform 1 0 696 0 1 570
box -8 -3 16 105
use FILL  FILL_4180
timestamp 1711653199
transform 1 0 688 0 1 570
box -8 -3 16 105
use FILL  FILL_4181
timestamp 1711653199
transform 1 0 680 0 1 570
box -8 -3 16 105
use FILL  FILL_4182
timestamp 1711653199
transform 1 0 640 0 1 570
box -8 -3 16 105
use FILL  FILL_4183
timestamp 1711653199
transform 1 0 632 0 1 570
box -8 -3 16 105
use FILL  FILL_4184
timestamp 1711653199
transform 1 0 608 0 1 570
box -8 -3 16 105
use FILL  FILL_4185
timestamp 1711653199
transform 1 0 600 0 1 570
box -8 -3 16 105
use FILL  FILL_4186
timestamp 1711653199
transform 1 0 592 0 1 570
box -8 -3 16 105
use FILL  FILL_4187
timestamp 1711653199
transform 1 0 552 0 1 570
box -8 -3 16 105
use FILL  FILL_4188
timestamp 1711653199
transform 1 0 544 0 1 570
box -8 -3 16 105
use FILL  FILL_4189
timestamp 1711653199
transform 1 0 504 0 1 570
box -8 -3 16 105
use FILL  FILL_4190
timestamp 1711653199
transform 1 0 496 0 1 570
box -8 -3 16 105
use FILL  FILL_4191
timestamp 1711653199
transform 1 0 488 0 1 570
box -8 -3 16 105
use FILL  FILL_4192
timestamp 1711653199
transform 1 0 480 0 1 570
box -8 -3 16 105
use FILL  FILL_4193
timestamp 1711653199
transform 1 0 440 0 1 570
box -8 -3 16 105
use FILL  FILL_4194
timestamp 1711653199
transform 1 0 432 0 1 570
box -8 -3 16 105
use FILL  FILL_4195
timestamp 1711653199
transform 1 0 424 0 1 570
box -8 -3 16 105
use FILL  FILL_4196
timestamp 1711653199
transform 1 0 376 0 1 570
box -8 -3 16 105
use FILL  FILL_4197
timestamp 1711653199
transform 1 0 368 0 1 570
box -8 -3 16 105
use FILL  FILL_4198
timestamp 1711653199
transform 1 0 360 0 1 570
box -8 -3 16 105
use FILL  FILL_4199
timestamp 1711653199
transform 1 0 352 0 1 570
box -8 -3 16 105
use FILL  FILL_4200
timestamp 1711653199
transform 1 0 344 0 1 570
box -8 -3 16 105
use FILL  FILL_4201
timestamp 1711653199
transform 1 0 336 0 1 570
box -8 -3 16 105
use FILL  FILL_4202
timestamp 1711653199
transform 1 0 280 0 1 570
box -8 -3 16 105
use FILL  FILL_4203
timestamp 1711653199
transform 1 0 272 0 1 570
box -8 -3 16 105
use FILL  FILL_4204
timestamp 1711653199
transform 1 0 264 0 1 570
box -8 -3 16 105
use FILL  FILL_4205
timestamp 1711653199
transform 1 0 256 0 1 570
box -8 -3 16 105
use FILL  FILL_4206
timestamp 1711653199
transform 1 0 208 0 1 570
box -8 -3 16 105
use FILL  FILL_4207
timestamp 1711653199
transform 1 0 200 0 1 570
box -8 -3 16 105
use FILL  FILL_4208
timestamp 1711653199
transform 1 0 192 0 1 570
box -8 -3 16 105
use FILL  FILL_4209
timestamp 1711653199
transform 1 0 184 0 1 570
box -8 -3 16 105
use FILL  FILL_4210
timestamp 1711653199
transform 1 0 176 0 1 570
box -8 -3 16 105
use FILL  FILL_4211
timestamp 1711653199
transform 1 0 128 0 1 570
box -8 -3 16 105
use FILL  FILL_4212
timestamp 1711653199
transform 1 0 120 0 1 570
box -8 -3 16 105
use FILL  FILL_4213
timestamp 1711653199
transform 1 0 112 0 1 570
box -8 -3 16 105
use FILL  FILL_4214
timestamp 1711653199
transform 1 0 80 0 1 570
box -8 -3 16 105
use FILL  FILL_4215
timestamp 1711653199
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_4216
timestamp 1711653199
transform 1 0 3392 0 -1 570
box -8 -3 16 105
use FILL  FILL_4217
timestamp 1711653199
transform 1 0 3384 0 -1 570
box -8 -3 16 105
use FILL  FILL_4218
timestamp 1711653199
transform 1 0 3344 0 -1 570
box -8 -3 16 105
use FILL  FILL_4219
timestamp 1711653199
transform 1 0 3336 0 -1 570
box -8 -3 16 105
use FILL  FILL_4220
timestamp 1711653199
transform 1 0 3328 0 -1 570
box -8 -3 16 105
use FILL  FILL_4221
timestamp 1711653199
transform 1 0 3320 0 -1 570
box -8 -3 16 105
use FILL  FILL_4222
timestamp 1711653199
transform 1 0 3296 0 -1 570
box -8 -3 16 105
use FILL  FILL_4223
timestamp 1711653199
transform 1 0 3264 0 -1 570
box -8 -3 16 105
use FILL  FILL_4224
timestamp 1711653199
transform 1 0 3256 0 -1 570
box -8 -3 16 105
use FILL  FILL_4225
timestamp 1711653199
transform 1 0 3248 0 -1 570
box -8 -3 16 105
use FILL  FILL_4226
timestamp 1711653199
transform 1 0 3240 0 -1 570
box -8 -3 16 105
use FILL  FILL_4227
timestamp 1711653199
transform 1 0 3232 0 -1 570
box -8 -3 16 105
use FILL  FILL_4228
timestamp 1711653199
transform 1 0 3184 0 -1 570
box -8 -3 16 105
use FILL  FILL_4229
timestamp 1711653199
transform 1 0 3176 0 -1 570
box -8 -3 16 105
use FILL  FILL_4230
timestamp 1711653199
transform 1 0 3168 0 -1 570
box -8 -3 16 105
use FILL  FILL_4231
timestamp 1711653199
transform 1 0 3160 0 -1 570
box -8 -3 16 105
use FILL  FILL_4232
timestamp 1711653199
transform 1 0 3120 0 -1 570
box -8 -3 16 105
use FILL  FILL_4233
timestamp 1711653199
transform 1 0 3112 0 -1 570
box -8 -3 16 105
use FILL  FILL_4234
timestamp 1711653199
transform 1 0 3104 0 -1 570
box -8 -3 16 105
use FILL  FILL_4235
timestamp 1711653199
transform 1 0 3096 0 -1 570
box -8 -3 16 105
use FILL  FILL_4236
timestamp 1711653199
transform 1 0 3064 0 -1 570
box -8 -3 16 105
use FILL  FILL_4237
timestamp 1711653199
transform 1 0 3032 0 -1 570
box -8 -3 16 105
use FILL  FILL_4238
timestamp 1711653199
transform 1 0 3024 0 -1 570
box -8 -3 16 105
use FILL  FILL_4239
timestamp 1711653199
transform 1 0 3016 0 -1 570
box -8 -3 16 105
use FILL  FILL_4240
timestamp 1711653199
transform 1 0 3008 0 -1 570
box -8 -3 16 105
use FILL  FILL_4241
timestamp 1711653199
transform 1 0 3000 0 -1 570
box -8 -3 16 105
use FILL  FILL_4242
timestamp 1711653199
transform 1 0 2992 0 -1 570
box -8 -3 16 105
use FILL  FILL_4243
timestamp 1711653199
transform 1 0 2968 0 -1 570
box -8 -3 16 105
use FILL  FILL_4244
timestamp 1711653199
transform 1 0 2944 0 -1 570
box -8 -3 16 105
use FILL  FILL_4245
timestamp 1711653199
transform 1 0 2936 0 -1 570
box -8 -3 16 105
use FILL  FILL_4246
timestamp 1711653199
transform 1 0 2904 0 -1 570
box -8 -3 16 105
use FILL  FILL_4247
timestamp 1711653199
transform 1 0 2896 0 -1 570
box -8 -3 16 105
use FILL  FILL_4248
timestamp 1711653199
transform 1 0 2888 0 -1 570
box -8 -3 16 105
use FILL  FILL_4249
timestamp 1711653199
transform 1 0 2880 0 -1 570
box -8 -3 16 105
use FILL  FILL_4250
timestamp 1711653199
transform 1 0 2872 0 -1 570
box -8 -3 16 105
use FILL  FILL_4251
timestamp 1711653199
transform 1 0 2816 0 -1 570
box -8 -3 16 105
use FILL  FILL_4252
timestamp 1711653199
transform 1 0 2808 0 -1 570
box -8 -3 16 105
use FILL  FILL_4253
timestamp 1711653199
transform 1 0 2800 0 -1 570
box -8 -3 16 105
use FILL  FILL_4254
timestamp 1711653199
transform 1 0 2792 0 -1 570
box -8 -3 16 105
use FILL  FILL_4255
timestamp 1711653199
transform 1 0 2784 0 -1 570
box -8 -3 16 105
use FILL  FILL_4256
timestamp 1711653199
transform 1 0 2776 0 -1 570
box -8 -3 16 105
use FILL  FILL_4257
timestamp 1711653199
transform 1 0 2768 0 -1 570
box -8 -3 16 105
use FILL  FILL_4258
timestamp 1711653199
transform 1 0 2712 0 -1 570
box -8 -3 16 105
use FILL  FILL_4259
timestamp 1711653199
transform 1 0 2704 0 -1 570
box -8 -3 16 105
use FILL  FILL_4260
timestamp 1711653199
transform 1 0 2696 0 -1 570
box -8 -3 16 105
use FILL  FILL_4261
timestamp 1711653199
transform 1 0 2688 0 -1 570
box -8 -3 16 105
use FILL  FILL_4262
timestamp 1711653199
transform 1 0 2656 0 -1 570
box -8 -3 16 105
use FILL  FILL_4263
timestamp 1711653199
transform 1 0 2648 0 -1 570
box -8 -3 16 105
use FILL  FILL_4264
timestamp 1711653199
transform 1 0 2600 0 -1 570
box -8 -3 16 105
use FILL  FILL_4265
timestamp 1711653199
transform 1 0 2592 0 -1 570
box -8 -3 16 105
use FILL  FILL_4266
timestamp 1711653199
transform 1 0 2584 0 -1 570
box -8 -3 16 105
use FILL  FILL_4267
timestamp 1711653199
transform 1 0 2576 0 -1 570
box -8 -3 16 105
use FILL  FILL_4268
timestamp 1711653199
transform 1 0 2528 0 -1 570
box -8 -3 16 105
use FILL  FILL_4269
timestamp 1711653199
transform 1 0 2520 0 -1 570
box -8 -3 16 105
use FILL  FILL_4270
timestamp 1711653199
transform 1 0 2512 0 -1 570
box -8 -3 16 105
use FILL  FILL_4271
timestamp 1711653199
transform 1 0 2472 0 -1 570
box -8 -3 16 105
use FILL  FILL_4272
timestamp 1711653199
transform 1 0 2464 0 -1 570
box -8 -3 16 105
use FILL  FILL_4273
timestamp 1711653199
transform 1 0 2456 0 -1 570
box -8 -3 16 105
use FILL  FILL_4274
timestamp 1711653199
transform 1 0 2448 0 -1 570
box -8 -3 16 105
use FILL  FILL_4275
timestamp 1711653199
transform 1 0 2440 0 -1 570
box -8 -3 16 105
use FILL  FILL_4276
timestamp 1711653199
transform 1 0 2432 0 -1 570
box -8 -3 16 105
use FILL  FILL_4277
timestamp 1711653199
transform 1 0 2384 0 -1 570
box -8 -3 16 105
use FILL  FILL_4278
timestamp 1711653199
transform 1 0 2376 0 -1 570
box -8 -3 16 105
use FILL  FILL_4279
timestamp 1711653199
transform 1 0 2368 0 -1 570
box -8 -3 16 105
use FILL  FILL_4280
timestamp 1711653199
transform 1 0 2360 0 -1 570
box -8 -3 16 105
use FILL  FILL_4281
timestamp 1711653199
transform 1 0 2336 0 -1 570
box -8 -3 16 105
use FILL  FILL_4282
timestamp 1711653199
transform 1 0 2328 0 -1 570
box -8 -3 16 105
use FILL  FILL_4283
timestamp 1711653199
transform 1 0 2320 0 -1 570
box -8 -3 16 105
use FILL  FILL_4284
timestamp 1711653199
transform 1 0 2312 0 -1 570
box -8 -3 16 105
use FILL  FILL_4285
timestamp 1711653199
transform 1 0 2304 0 -1 570
box -8 -3 16 105
use FILL  FILL_4286
timestamp 1711653199
transform 1 0 2256 0 -1 570
box -8 -3 16 105
use FILL  FILL_4287
timestamp 1711653199
transform 1 0 2248 0 -1 570
box -8 -3 16 105
use FILL  FILL_4288
timestamp 1711653199
transform 1 0 2240 0 -1 570
box -8 -3 16 105
use FILL  FILL_4289
timestamp 1711653199
transform 1 0 2232 0 -1 570
box -8 -3 16 105
use FILL  FILL_4290
timestamp 1711653199
transform 1 0 2200 0 -1 570
box -8 -3 16 105
use FILL  FILL_4291
timestamp 1711653199
transform 1 0 2192 0 -1 570
box -8 -3 16 105
use FILL  FILL_4292
timestamp 1711653199
transform 1 0 2184 0 -1 570
box -8 -3 16 105
use FILL  FILL_4293
timestamp 1711653199
transform 1 0 2176 0 -1 570
box -8 -3 16 105
use FILL  FILL_4294
timestamp 1711653199
transform 1 0 2168 0 -1 570
box -8 -3 16 105
use FILL  FILL_4295
timestamp 1711653199
transform 1 0 2160 0 -1 570
box -8 -3 16 105
use FILL  FILL_4296
timestamp 1711653199
transform 1 0 2112 0 -1 570
box -8 -3 16 105
use FILL  FILL_4297
timestamp 1711653199
transform 1 0 2104 0 -1 570
box -8 -3 16 105
use FILL  FILL_4298
timestamp 1711653199
transform 1 0 2096 0 -1 570
box -8 -3 16 105
use FILL  FILL_4299
timestamp 1711653199
transform 1 0 2088 0 -1 570
box -8 -3 16 105
use FILL  FILL_4300
timestamp 1711653199
transform 1 0 2080 0 -1 570
box -8 -3 16 105
use FILL  FILL_4301
timestamp 1711653199
transform 1 0 2048 0 -1 570
box -8 -3 16 105
use FILL  FILL_4302
timestamp 1711653199
transform 1 0 2040 0 -1 570
box -8 -3 16 105
use FILL  FILL_4303
timestamp 1711653199
transform 1 0 2032 0 -1 570
box -8 -3 16 105
use FILL  FILL_4304
timestamp 1711653199
transform 1 0 1992 0 -1 570
box -8 -3 16 105
use FILL  FILL_4305
timestamp 1711653199
transform 1 0 1984 0 -1 570
box -8 -3 16 105
use FILL  FILL_4306
timestamp 1711653199
transform 1 0 1976 0 -1 570
box -8 -3 16 105
use FILL  FILL_4307
timestamp 1711653199
transform 1 0 1968 0 -1 570
box -8 -3 16 105
use FILL  FILL_4308
timestamp 1711653199
transform 1 0 1960 0 -1 570
box -8 -3 16 105
use FILL  FILL_4309
timestamp 1711653199
transform 1 0 1952 0 -1 570
box -8 -3 16 105
use FILL  FILL_4310
timestamp 1711653199
transform 1 0 1944 0 -1 570
box -8 -3 16 105
use FILL  FILL_4311
timestamp 1711653199
transform 1 0 1896 0 -1 570
box -8 -3 16 105
use FILL  FILL_4312
timestamp 1711653199
transform 1 0 1888 0 -1 570
box -8 -3 16 105
use FILL  FILL_4313
timestamp 1711653199
transform 1 0 1880 0 -1 570
box -8 -3 16 105
use FILL  FILL_4314
timestamp 1711653199
transform 1 0 1872 0 -1 570
box -8 -3 16 105
use FILL  FILL_4315
timestamp 1711653199
transform 1 0 1864 0 -1 570
box -8 -3 16 105
use FILL  FILL_4316
timestamp 1711653199
transform 1 0 1832 0 -1 570
box -8 -3 16 105
use FILL  FILL_4317
timestamp 1711653199
transform 1 0 1824 0 -1 570
box -8 -3 16 105
use FILL  FILL_4318
timestamp 1711653199
transform 1 0 1816 0 -1 570
box -8 -3 16 105
use FILL  FILL_4319
timestamp 1711653199
transform 1 0 1808 0 -1 570
box -8 -3 16 105
use FILL  FILL_4320
timestamp 1711653199
transform 1 0 1776 0 -1 570
box -8 -3 16 105
use FILL  FILL_4321
timestamp 1711653199
transform 1 0 1768 0 -1 570
box -8 -3 16 105
use FILL  FILL_4322
timestamp 1711653199
transform 1 0 1760 0 -1 570
box -8 -3 16 105
use FILL  FILL_4323
timestamp 1711653199
transform 1 0 1752 0 -1 570
box -8 -3 16 105
use FILL  FILL_4324
timestamp 1711653199
transform 1 0 1744 0 -1 570
box -8 -3 16 105
use FILL  FILL_4325
timestamp 1711653199
transform 1 0 1736 0 -1 570
box -8 -3 16 105
use FILL  FILL_4326
timestamp 1711653199
transform 1 0 1688 0 -1 570
box -8 -3 16 105
use FILL  FILL_4327
timestamp 1711653199
transform 1 0 1680 0 -1 570
box -8 -3 16 105
use FILL  FILL_4328
timestamp 1711653199
transform 1 0 1672 0 -1 570
box -8 -3 16 105
use FILL  FILL_4329
timestamp 1711653199
transform 1 0 1664 0 -1 570
box -8 -3 16 105
use FILL  FILL_4330
timestamp 1711653199
transform 1 0 1656 0 -1 570
box -8 -3 16 105
use FILL  FILL_4331
timestamp 1711653199
transform 1 0 1648 0 -1 570
box -8 -3 16 105
use FILL  FILL_4332
timestamp 1711653199
transform 1 0 1640 0 -1 570
box -8 -3 16 105
use FILL  FILL_4333
timestamp 1711653199
transform 1 0 1600 0 -1 570
box -8 -3 16 105
use FILL  FILL_4334
timestamp 1711653199
transform 1 0 1592 0 -1 570
box -8 -3 16 105
use FILL  FILL_4335
timestamp 1711653199
transform 1 0 1584 0 -1 570
box -8 -3 16 105
use FILL  FILL_4336
timestamp 1711653199
transform 1 0 1576 0 -1 570
box -8 -3 16 105
use FILL  FILL_4337
timestamp 1711653199
transform 1 0 1568 0 -1 570
box -8 -3 16 105
use FILL  FILL_4338
timestamp 1711653199
transform 1 0 1528 0 -1 570
box -8 -3 16 105
use FILL  FILL_4339
timestamp 1711653199
transform 1 0 1520 0 -1 570
box -8 -3 16 105
use FILL  FILL_4340
timestamp 1711653199
transform 1 0 1512 0 -1 570
box -8 -3 16 105
use FILL  FILL_4341
timestamp 1711653199
transform 1 0 1504 0 -1 570
box -8 -3 16 105
use FILL  FILL_4342
timestamp 1711653199
transform 1 0 1496 0 -1 570
box -8 -3 16 105
use FILL  FILL_4343
timestamp 1711653199
transform 1 0 1488 0 -1 570
box -8 -3 16 105
use FILL  FILL_4344
timestamp 1711653199
transform 1 0 1448 0 -1 570
box -8 -3 16 105
use FILL  FILL_4345
timestamp 1711653199
transform 1 0 1440 0 -1 570
box -8 -3 16 105
use FILL  FILL_4346
timestamp 1711653199
transform 1 0 1432 0 -1 570
box -8 -3 16 105
use FILL  FILL_4347
timestamp 1711653199
transform 1 0 1424 0 -1 570
box -8 -3 16 105
use FILL  FILL_4348
timestamp 1711653199
transform 1 0 1416 0 -1 570
box -8 -3 16 105
use FILL  FILL_4349
timestamp 1711653199
transform 1 0 1384 0 -1 570
box -8 -3 16 105
use FILL  FILL_4350
timestamp 1711653199
transform 1 0 1376 0 -1 570
box -8 -3 16 105
use FILL  FILL_4351
timestamp 1711653199
transform 1 0 1368 0 -1 570
box -8 -3 16 105
use FILL  FILL_4352
timestamp 1711653199
transform 1 0 1360 0 -1 570
box -8 -3 16 105
use FILL  FILL_4353
timestamp 1711653199
transform 1 0 1352 0 -1 570
box -8 -3 16 105
use FILL  FILL_4354
timestamp 1711653199
transform 1 0 1312 0 -1 570
box -8 -3 16 105
use FILL  FILL_4355
timestamp 1711653199
transform 1 0 1304 0 -1 570
box -8 -3 16 105
use FILL  FILL_4356
timestamp 1711653199
transform 1 0 1296 0 -1 570
box -8 -3 16 105
use FILL  FILL_4357
timestamp 1711653199
transform 1 0 1288 0 -1 570
box -8 -3 16 105
use FILL  FILL_4358
timestamp 1711653199
transform 1 0 1280 0 -1 570
box -8 -3 16 105
use FILL  FILL_4359
timestamp 1711653199
transform 1 0 1272 0 -1 570
box -8 -3 16 105
use FILL  FILL_4360
timestamp 1711653199
transform 1 0 1264 0 -1 570
box -8 -3 16 105
use FILL  FILL_4361
timestamp 1711653199
transform 1 0 1224 0 -1 570
box -8 -3 16 105
use FILL  FILL_4362
timestamp 1711653199
transform 1 0 1216 0 -1 570
box -8 -3 16 105
use FILL  FILL_4363
timestamp 1711653199
transform 1 0 1208 0 -1 570
box -8 -3 16 105
use FILL  FILL_4364
timestamp 1711653199
transform 1 0 1200 0 -1 570
box -8 -3 16 105
use FILL  FILL_4365
timestamp 1711653199
transform 1 0 1176 0 -1 570
box -8 -3 16 105
use FILL  FILL_4366
timestamp 1711653199
transform 1 0 1168 0 -1 570
box -8 -3 16 105
use FILL  FILL_4367
timestamp 1711653199
transform 1 0 1160 0 -1 570
box -8 -3 16 105
use FILL  FILL_4368
timestamp 1711653199
transform 1 0 1152 0 -1 570
box -8 -3 16 105
use FILL  FILL_4369
timestamp 1711653199
transform 1 0 1112 0 -1 570
box -8 -3 16 105
use FILL  FILL_4370
timestamp 1711653199
transform 1 0 1104 0 -1 570
box -8 -3 16 105
use FILL  FILL_4371
timestamp 1711653199
transform 1 0 1096 0 -1 570
box -8 -3 16 105
use FILL  FILL_4372
timestamp 1711653199
transform 1 0 1088 0 -1 570
box -8 -3 16 105
use FILL  FILL_4373
timestamp 1711653199
transform 1 0 1080 0 -1 570
box -8 -3 16 105
use FILL  FILL_4374
timestamp 1711653199
transform 1 0 1040 0 -1 570
box -8 -3 16 105
use FILL  FILL_4375
timestamp 1711653199
transform 1 0 1032 0 -1 570
box -8 -3 16 105
use FILL  FILL_4376
timestamp 1711653199
transform 1 0 1024 0 -1 570
box -8 -3 16 105
use FILL  FILL_4377
timestamp 1711653199
transform 1 0 1016 0 -1 570
box -8 -3 16 105
use FILL  FILL_4378
timestamp 1711653199
transform 1 0 1008 0 -1 570
box -8 -3 16 105
use FILL  FILL_4379
timestamp 1711653199
transform 1 0 1000 0 -1 570
box -8 -3 16 105
use FILL  FILL_4380
timestamp 1711653199
transform 1 0 960 0 -1 570
box -8 -3 16 105
use FILL  FILL_4381
timestamp 1711653199
transform 1 0 952 0 -1 570
box -8 -3 16 105
use FILL  FILL_4382
timestamp 1711653199
transform 1 0 928 0 -1 570
box -8 -3 16 105
use FILL  FILL_4383
timestamp 1711653199
transform 1 0 920 0 -1 570
box -8 -3 16 105
use FILL  FILL_4384
timestamp 1711653199
transform 1 0 912 0 -1 570
box -8 -3 16 105
use FILL  FILL_4385
timestamp 1711653199
transform 1 0 904 0 -1 570
box -8 -3 16 105
use FILL  FILL_4386
timestamp 1711653199
transform 1 0 896 0 -1 570
box -8 -3 16 105
use FILL  FILL_4387
timestamp 1711653199
transform 1 0 888 0 -1 570
box -8 -3 16 105
use FILL  FILL_4388
timestamp 1711653199
transform 1 0 864 0 -1 570
box -8 -3 16 105
use FILL  FILL_4389
timestamp 1711653199
transform 1 0 856 0 -1 570
box -8 -3 16 105
use FILL  FILL_4390
timestamp 1711653199
transform 1 0 808 0 -1 570
box -8 -3 16 105
use FILL  FILL_4391
timestamp 1711653199
transform 1 0 800 0 -1 570
box -8 -3 16 105
use FILL  FILL_4392
timestamp 1711653199
transform 1 0 792 0 -1 570
box -8 -3 16 105
use FILL  FILL_4393
timestamp 1711653199
transform 1 0 784 0 -1 570
box -8 -3 16 105
use FILL  FILL_4394
timestamp 1711653199
transform 1 0 776 0 -1 570
box -8 -3 16 105
use FILL  FILL_4395
timestamp 1711653199
transform 1 0 768 0 -1 570
box -8 -3 16 105
use FILL  FILL_4396
timestamp 1711653199
transform 1 0 760 0 -1 570
box -8 -3 16 105
use FILL  FILL_4397
timestamp 1711653199
transform 1 0 688 0 -1 570
box -8 -3 16 105
use FILL  FILL_4398
timestamp 1711653199
transform 1 0 680 0 -1 570
box -8 -3 16 105
use FILL  FILL_4399
timestamp 1711653199
transform 1 0 672 0 -1 570
box -8 -3 16 105
use FILL  FILL_4400
timestamp 1711653199
transform 1 0 664 0 -1 570
box -8 -3 16 105
use FILL  FILL_4401
timestamp 1711653199
transform 1 0 656 0 -1 570
box -8 -3 16 105
use FILL  FILL_4402
timestamp 1711653199
transform 1 0 648 0 -1 570
box -8 -3 16 105
use FILL  FILL_4403
timestamp 1711653199
transform 1 0 640 0 -1 570
box -8 -3 16 105
use FILL  FILL_4404
timestamp 1711653199
transform 1 0 584 0 -1 570
box -8 -3 16 105
use FILL  FILL_4405
timestamp 1711653199
transform 1 0 576 0 -1 570
box -8 -3 16 105
use FILL  FILL_4406
timestamp 1711653199
transform 1 0 568 0 -1 570
box -8 -3 16 105
use FILL  FILL_4407
timestamp 1711653199
transform 1 0 560 0 -1 570
box -8 -3 16 105
use FILL  FILL_4408
timestamp 1711653199
transform 1 0 552 0 -1 570
box -8 -3 16 105
use FILL  FILL_4409
timestamp 1711653199
transform 1 0 544 0 -1 570
box -8 -3 16 105
use FILL  FILL_4410
timestamp 1711653199
transform 1 0 536 0 -1 570
box -8 -3 16 105
use FILL  FILL_4411
timestamp 1711653199
transform 1 0 480 0 -1 570
box -8 -3 16 105
use FILL  FILL_4412
timestamp 1711653199
transform 1 0 472 0 -1 570
box -8 -3 16 105
use FILL  FILL_4413
timestamp 1711653199
transform 1 0 464 0 -1 570
box -8 -3 16 105
use FILL  FILL_4414
timestamp 1711653199
transform 1 0 456 0 -1 570
box -8 -3 16 105
use FILL  FILL_4415
timestamp 1711653199
transform 1 0 448 0 -1 570
box -8 -3 16 105
use FILL  FILL_4416
timestamp 1711653199
transform 1 0 440 0 -1 570
box -8 -3 16 105
use FILL  FILL_4417
timestamp 1711653199
transform 1 0 432 0 -1 570
box -8 -3 16 105
use FILL  FILL_4418
timestamp 1711653199
transform 1 0 424 0 -1 570
box -8 -3 16 105
use FILL  FILL_4419
timestamp 1711653199
transform 1 0 376 0 -1 570
box -8 -3 16 105
use FILL  FILL_4420
timestamp 1711653199
transform 1 0 368 0 -1 570
box -8 -3 16 105
use FILL  FILL_4421
timestamp 1711653199
transform 1 0 360 0 -1 570
box -8 -3 16 105
use FILL  FILL_4422
timestamp 1711653199
transform 1 0 352 0 -1 570
box -8 -3 16 105
use FILL  FILL_4423
timestamp 1711653199
transform 1 0 344 0 -1 570
box -8 -3 16 105
use FILL  FILL_4424
timestamp 1711653199
transform 1 0 336 0 -1 570
box -8 -3 16 105
use FILL  FILL_4425
timestamp 1711653199
transform 1 0 328 0 -1 570
box -8 -3 16 105
use FILL  FILL_4426
timestamp 1711653199
transform 1 0 280 0 -1 570
box -8 -3 16 105
use FILL  FILL_4427
timestamp 1711653199
transform 1 0 272 0 -1 570
box -8 -3 16 105
use FILL  FILL_4428
timestamp 1711653199
transform 1 0 264 0 -1 570
box -8 -3 16 105
use FILL  FILL_4429
timestamp 1711653199
transform 1 0 256 0 -1 570
box -8 -3 16 105
use FILL  FILL_4430
timestamp 1711653199
transform 1 0 248 0 -1 570
box -8 -3 16 105
use FILL  FILL_4431
timestamp 1711653199
transform 1 0 240 0 -1 570
box -8 -3 16 105
use FILL  FILL_4432
timestamp 1711653199
transform 1 0 232 0 -1 570
box -8 -3 16 105
use FILL  FILL_4433
timestamp 1711653199
transform 1 0 184 0 -1 570
box -8 -3 16 105
use FILL  FILL_4434
timestamp 1711653199
transform 1 0 176 0 -1 570
box -8 -3 16 105
use FILL  FILL_4435
timestamp 1711653199
transform 1 0 168 0 -1 570
box -8 -3 16 105
use FILL  FILL_4436
timestamp 1711653199
transform 1 0 160 0 -1 570
box -8 -3 16 105
use FILL  FILL_4437
timestamp 1711653199
transform 1 0 152 0 -1 570
box -8 -3 16 105
use FILL  FILL_4438
timestamp 1711653199
transform 1 0 120 0 -1 570
box -8 -3 16 105
use FILL  FILL_4439
timestamp 1711653199
transform 1 0 112 0 -1 570
box -8 -3 16 105
use FILL  FILL_4440
timestamp 1711653199
transform 1 0 104 0 -1 570
box -8 -3 16 105
use FILL  FILL_4441
timestamp 1711653199
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_4442
timestamp 1711653199
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_4443
timestamp 1711653199
transform 1 0 3392 0 1 370
box -8 -3 16 105
use FILL  FILL_4444
timestamp 1711653199
transform 1 0 3384 0 1 370
box -8 -3 16 105
use FILL  FILL_4445
timestamp 1711653199
transform 1 0 3376 0 1 370
box -8 -3 16 105
use FILL  FILL_4446
timestamp 1711653199
transform 1 0 3336 0 1 370
box -8 -3 16 105
use FILL  FILL_4447
timestamp 1711653199
transform 1 0 3304 0 1 370
box -8 -3 16 105
use FILL  FILL_4448
timestamp 1711653199
transform 1 0 3296 0 1 370
box -8 -3 16 105
use FILL  FILL_4449
timestamp 1711653199
transform 1 0 3288 0 1 370
box -8 -3 16 105
use FILL  FILL_4450
timestamp 1711653199
transform 1 0 3280 0 1 370
box -8 -3 16 105
use FILL  FILL_4451
timestamp 1711653199
transform 1 0 3248 0 1 370
box -8 -3 16 105
use FILL  FILL_4452
timestamp 1711653199
transform 1 0 3240 0 1 370
box -8 -3 16 105
use FILL  FILL_4453
timestamp 1711653199
transform 1 0 3232 0 1 370
box -8 -3 16 105
use FILL  FILL_4454
timestamp 1711653199
transform 1 0 3184 0 1 370
box -8 -3 16 105
use FILL  FILL_4455
timestamp 1711653199
transform 1 0 3176 0 1 370
box -8 -3 16 105
use FILL  FILL_4456
timestamp 1711653199
transform 1 0 3168 0 1 370
box -8 -3 16 105
use FILL  FILL_4457
timestamp 1711653199
transform 1 0 3160 0 1 370
box -8 -3 16 105
use FILL  FILL_4458
timestamp 1711653199
transform 1 0 3152 0 1 370
box -8 -3 16 105
use FILL  FILL_4459
timestamp 1711653199
transform 1 0 3144 0 1 370
box -8 -3 16 105
use FILL  FILL_4460
timestamp 1711653199
transform 1 0 3096 0 1 370
box -8 -3 16 105
use FILL  FILL_4461
timestamp 1711653199
transform 1 0 3088 0 1 370
box -8 -3 16 105
use FILL  FILL_4462
timestamp 1711653199
transform 1 0 3080 0 1 370
box -8 -3 16 105
use FILL  FILL_4463
timestamp 1711653199
transform 1 0 3072 0 1 370
box -8 -3 16 105
use FILL  FILL_4464
timestamp 1711653199
transform 1 0 3016 0 1 370
box -8 -3 16 105
use FILL  FILL_4465
timestamp 1711653199
transform 1 0 3008 0 1 370
box -8 -3 16 105
use FILL  FILL_4466
timestamp 1711653199
transform 1 0 3000 0 1 370
box -8 -3 16 105
use FILL  FILL_4467
timestamp 1711653199
transform 1 0 2992 0 1 370
box -8 -3 16 105
use FILL  FILL_4468
timestamp 1711653199
transform 1 0 2984 0 1 370
box -8 -3 16 105
use FILL  FILL_4469
timestamp 1711653199
transform 1 0 2976 0 1 370
box -8 -3 16 105
use FILL  FILL_4470
timestamp 1711653199
transform 1 0 2912 0 1 370
box -8 -3 16 105
use FILL  FILL_4471
timestamp 1711653199
transform 1 0 2904 0 1 370
box -8 -3 16 105
use FILL  FILL_4472
timestamp 1711653199
transform 1 0 2896 0 1 370
box -8 -3 16 105
use FILL  FILL_4473
timestamp 1711653199
transform 1 0 2888 0 1 370
box -8 -3 16 105
use FILL  FILL_4474
timestamp 1711653199
transform 1 0 2880 0 1 370
box -8 -3 16 105
use FILL  FILL_4475
timestamp 1711653199
transform 1 0 2872 0 1 370
box -8 -3 16 105
use FILL  FILL_4476
timestamp 1711653199
transform 1 0 2824 0 1 370
box -8 -3 16 105
use FILL  FILL_4477
timestamp 1711653199
transform 1 0 2816 0 1 370
box -8 -3 16 105
use FILL  FILL_4478
timestamp 1711653199
transform 1 0 2768 0 1 370
box -8 -3 16 105
use FILL  FILL_4479
timestamp 1711653199
transform 1 0 2760 0 1 370
box -8 -3 16 105
use FILL  FILL_4480
timestamp 1711653199
transform 1 0 2752 0 1 370
box -8 -3 16 105
use FILL  FILL_4481
timestamp 1711653199
transform 1 0 2744 0 1 370
box -8 -3 16 105
use FILL  FILL_4482
timestamp 1711653199
transform 1 0 2736 0 1 370
box -8 -3 16 105
use FILL  FILL_4483
timestamp 1711653199
transform 1 0 2672 0 1 370
box -8 -3 16 105
use FILL  FILL_4484
timestamp 1711653199
transform 1 0 2664 0 1 370
box -8 -3 16 105
use FILL  FILL_4485
timestamp 1711653199
transform 1 0 2656 0 1 370
box -8 -3 16 105
use FILL  FILL_4486
timestamp 1711653199
transform 1 0 2648 0 1 370
box -8 -3 16 105
use FILL  FILL_4487
timestamp 1711653199
transform 1 0 2600 0 1 370
box -8 -3 16 105
use FILL  FILL_4488
timestamp 1711653199
transform 1 0 2592 0 1 370
box -8 -3 16 105
use FILL  FILL_4489
timestamp 1711653199
transform 1 0 2584 0 1 370
box -8 -3 16 105
use FILL  FILL_4490
timestamp 1711653199
transform 1 0 2576 0 1 370
box -8 -3 16 105
use FILL  FILL_4491
timestamp 1711653199
transform 1 0 2568 0 1 370
box -8 -3 16 105
use FILL  FILL_4492
timestamp 1711653199
transform 1 0 2536 0 1 370
box -8 -3 16 105
use FILL  FILL_4493
timestamp 1711653199
transform 1 0 2528 0 1 370
box -8 -3 16 105
use FILL  FILL_4494
timestamp 1711653199
transform 1 0 2520 0 1 370
box -8 -3 16 105
use FILL  FILL_4495
timestamp 1711653199
transform 1 0 2512 0 1 370
box -8 -3 16 105
use FILL  FILL_4496
timestamp 1711653199
transform 1 0 2464 0 1 370
box -8 -3 16 105
use FILL  FILL_4497
timestamp 1711653199
transform 1 0 2456 0 1 370
box -8 -3 16 105
use FILL  FILL_4498
timestamp 1711653199
transform 1 0 2448 0 1 370
box -8 -3 16 105
use FILL  FILL_4499
timestamp 1711653199
transform 1 0 2440 0 1 370
box -8 -3 16 105
use FILL  FILL_4500
timestamp 1711653199
transform 1 0 2432 0 1 370
box -8 -3 16 105
use FILL  FILL_4501
timestamp 1711653199
transform 1 0 2392 0 1 370
box -8 -3 16 105
use FILL  FILL_4502
timestamp 1711653199
transform 1 0 2384 0 1 370
box -8 -3 16 105
use FILL  FILL_4503
timestamp 1711653199
transform 1 0 2376 0 1 370
box -8 -3 16 105
use FILL  FILL_4504
timestamp 1711653199
transform 1 0 2368 0 1 370
box -8 -3 16 105
use FILL  FILL_4505
timestamp 1711653199
transform 1 0 2360 0 1 370
box -8 -3 16 105
use FILL  FILL_4506
timestamp 1711653199
transform 1 0 2320 0 1 370
box -8 -3 16 105
use FILL  FILL_4507
timestamp 1711653199
transform 1 0 2312 0 1 370
box -8 -3 16 105
use FILL  FILL_4508
timestamp 1711653199
transform 1 0 2304 0 1 370
box -8 -3 16 105
use FILL  FILL_4509
timestamp 1711653199
transform 1 0 2296 0 1 370
box -8 -3 16 105
use FILL  FILL_4510
timestamp 1711653199
transform 1 0 2288 0 1 370
box -8 -3 16 105
use FILL  FILL_4511
timestamp 1711653199
transform 1 0 2240 0 1 370
box -8 -3 16 105
use FILL  FILL_4512
timestamp 1711653199
transform 1 0 2232 0 1 370
box -8 -3 16 105
use FILL  FILL_4513
timestamp 1711653199
transform 1 0 2224 0 1 370
box -8 -3 16 105
use FILL  FILL_4514
timestamp 1711653199
transform 1 0 2216 0 1 370
box -8 -3 16 105
use FILL  FILL_4515
timestamp 1711653199
transform 1 0 2208 0 1 370
box -8 -3 16 105
use FILL  FILL_4516
timestamp 1711653199
transform 1 0 2200 0 1 370
box -8 -3 16 105
use FILL  FILL_4517
timestamp 1711653199
transform 1 0 2160 0 1 370
box -8 -3 16 105
use FILL  FILL_4518
timestamp 1711653199
transform 1 0 2152 0 1 370
box -8 -3 16 105
use FILL  FILL_4519
timestamp 1711653199
transform 1 0 2144 0 1 370
box -8 -3 16 105
use FILL  FILL_4520
timestamp 1711653199
transform 1 0 2136 0 1 370
box -8 -3 16 105
use FILL  FILL_4521
timestamp 1711653199
transform 1 0 2096 0 1 370
box -8 -3 16 105
use FILL  FILL_4522
timestamp 1711653199
transform 1 0 2088 0 1 370
box -8 -3 16 105
use FILL  FILL_4523
timestamp 1711653199
transform 1 0 2080 0 1 370
box -8 -3 16 105
use FILL  FILL_4524
timestamp 1711653199
transform 1 0 2072 0 1 370
box -8 -3 16 105
use FILL  FILL_4525
timestamp 1711653199
transform 1 0 2064 0 1 370
box -8 -3 16 105
use FILL  FILL_4526
timestamp 1711653199
transform 1 0 1992 0 1 370
box -8 -3 16 105
use FILL  FILL_4527
timestamp 1711653199
transform 1 0 1984 0 1 370
box -8 -3 16 105
use FILL  FILL_4528
timestamp 1711653199
transform 1 0 1976 0 1 370
box -8 -3 16 105
use FILL  FILL_4529
timestamp 1711653199
transform 1 0 1968 0 1 370
box -8 -3 16 105
use FILL  FILL_4530
timestamp 1711653199
transform 1 0 1960 0 1 370
box -8 -3 16 105
use FILL  FILL_4531
timestamp 1711653199
transform 1 0 1936 0 1 370
box -8 -3 16 105
use FILL  FILL_4532
timestamp 1711653199
transform 1 0 1904 0 1 370
box -8 -3 16 105
use FILL  FILL_4533
timestamp 1711653199
transform 1 0 1896 0 1 370
box -8 -3 16 105
use FILL  FILL_4534
timestamp 1711653199
transform 1 0 1888 0 1 370
box -8 -3 16 105
use FILL  FILL_4535
timestamp 1711653199
transform 1 0 1880 0 1 370
box -8 -3 16 105
use FILL  FILL_4536
timestamp 1711653199
transform 1 0 1872 0 1 370
box -8 -3 16 105
use FILL  FILL_4537
timestamp 1711653199
transform 1 0 1848 0 1 370
box -8 -3 16 105
use FILL  FILL_4538
timestamp 1711653199
transform 1 0 1840 0 1 370
box -8 -3 16 105
use FILL  FILL_4539
timestamp 1711653199
transform 1 0 1832 0 1 370
box -8 -3 16 105
use FILL  FILL_4540
timestamp 1711653199
transform 1 0 1800 0 1 370
box -8 -3 16 105
use FILL  FILL_4541
timestamp 1711653199
transform 1 0 1792 0 1 370
box -8 -3 16 105
use FILL  FILL_4542
timestamp 1711653199
transform 1 0 1784 0 1 370
box -8 -3 16 105
use FILL  FILL_4543
timestamp 1711653199
transform 1 0 1776 0 1 370
box -8 -3 16 105
use FILL  FILL_4544
timestamp 1711653199
transform 1 0 1768 0 1 370
box -8 -3 16 105
use FILL  FILL_4545
timestamp 1711653199
transform 1 0 1728 0 1 370
box -8 -3 16 105
use FILL  FILL_4546
timestamp 1711653199
transform 1 0 1720 0 1 370
box -8 -3 16 105
use FILL  FILL_4547
timestamp 1711653199
transform 1 0 1712 0 1 370
box -8 -3 16 105
use FILL  FILL_4548
timestamp 1711653199
transform 1 0 1704 0 1 370
box -8 -3 16 105
use FILL  FILL_4549
timestamp 1711653199
transform 1 0 1696 0 1 370
box -8 -3 16 105
use FILL  FILL_4550
timestamp 1711653199
transform 1 0 1664 0 1 370
box -8 -3 16 105
use FILL  FILL_4551
timestamp 1711653199
transform 1 0 1656 0 1 370
box -8 -3 16 105
use FILL  FILL_4552
timestamp 1711653199
transform 1 0 1648 0 1 370
box -8 -3 16 105
use FILL  FILL_4553
timestamp 1711653199
transform 1 0 1640 0 1 370
box -8 -3 16 105
use FILL  FILL_4554
timestamp 1711653199
transform 1 0 1632 0 1 370
box -8 -3 16 105
use FILL  FILL_4555
timestamp 1711653199
transform 1 0 1600 0 1 370
box -8 -3 16 105
use FILL  FILL_4556
timestamp 1711653199
transform 1 0 1592 0 1 370
box -8 -3 16 105
use FILL  FILL_4557
timestamp 1711653199
transform 1 0 1584 0 1 370
box -8 -3 16 105
use FILL  FILL_4558
timestamp 1711653199
transform 1 0 1576 0 1 370
box -8 -3 16 105
use FILL  FILL_4559
timestamp 1711653199
transform 1 0 1568 0 1 370
box -8 -3 16 105
use FILL  FILL_4560
timestamp 1711653199
transform 1 0 1528 0 1 370
box -8 -3 16 105
use FILL  FILL_4561
timestamp 1711653199
transform 1 0 1520 0 1 370
box -8 -3 16 105
use FILL  FILL_4562
timestamp 1711653199
transform 1 0 1512 0 1 370
box -8 -3 16 105
use FILL  FILL_4563
timestamp 1711653199
transform 1 0 1504 0 1 370
box -8 -3 16 105
use FILL  FILL_4564
timestamp 1711653199
transform 1 0 1496 0 1 370
box -8 -3 16 105
use FILL  FILL_4565
timestamp 1711653199
transform 1 0 1456 0 1 370
box -8 -3 16 105
use FILL  FILL_4566
timestamp 1711653199
transform 1 0 1448 0 1 370
box -8 -3 16 105
use FILL  FILL_4567
timestamp 1711653199
transform 1 0 1440 0 1 370
box -8 -3 16 105
use FILL  FILL_4568
timestamp 1711653199
transform 1 0 1432 0 1 370
box -8 -3 16 105
use FILL  FILL_4569
timestamp 1711653199
transform 1 0 1424 0 1 370
box -8 -3 16 105
use FILL  FILL_4570
timestamp 1711653199
transform 1 0 1384 0 1 370
box -8 -3 16 105
use FILL  FILL_4571
timestamp 1711653199
transform 1 0 1376 0 1 370
box -8 -3 16 105
use FILL  FILL_4572
timestamp 1711653199
transform 1 0 1368 0 1 370
box -8 -3 16 105
use FILL  FILL_4573
timestamp 1711653199
transform 1 0 1336 0 1 370
box -8 -3 16 105
use FILL  FILL_4574
timestamp 1711653199
transform 1 0 1312 0 1 370
box -8 -3 16 105
use FILL  FILL_4575
timestamp 1711653199
transform 1 0 1304 0 1 370
box -8 -3 16 105
use FILL  FILL_4576
timestamp 1711653199
transform 1 0 1296 0 1 370
box -8 -3 16 105
use FILL  FILL_4577
timestamp 1711653199
transform 1 0 1288 0 1 370
box -8 -3 16 105
use FILL  FILL_4578
timestamp 1711653199
transform 1 0 1280 0 1 370
box -8 -3 16 105
use FILL  FILL_4579
timestamp 1711653199
transform 1 0 1272 0 1 370
box -8 -3 16 105
use FILL  FILL_4580
timestamp 1711653199
transform 1 0 1224 0 1 370
box -8 -3 16 105
use FILL  FILL_4581
timestamp 1711653199
transform 1 0 1216 0 1 370
box -8 -3 16 105
use FILL  FILL_4582
timestamp 1711653199
transform 1 0 1208 0 1 370
box -8 -3 16 105
use FILL  FILL_4583
timestamp 1711653199
transform 1 0 1200 0 1 370
box -8 -3 16 105
use FILL  FILL_4584
timestamp 1711653199
transform 1 0 1192 0 1 370
box -8 -3 16 105
use FILL  FILL_4585
timestamp 1711653199
transform 1 0 1152 0 1 370
box -8 -3 16 105
use FILL  FILL_4586
timestamp 1711653199
transform 1 0 1144 0 1 370
box -8 -3 16 105
use FILL  FILL_4587
timestamp 1711653199
transform 1 0 1104 0 1 370
box -8 -3 16 105
use FILL  FILL_4588
timestamp 1711653199
transform 1 0 1096 0 1 370
box -8 -3 16 105
use FILL  FILL_4589
timestamp 1711653199
transform 1 0 1088 0 1 370
box -8 -3 16 105
use FILL  FILL_4590
timestamp 1711653199
transform 1 0 1048 0 1 370
box -8 -3 16 105
use FILL  FILL_4591
timestamp 1711653199
transform 1 0 1040 0 1 370
box -8 -3 16 105
use FILL  FILL_4592
timestamp 1711653199
transform 1 0 1032 0 1 370
box -8 -3 16 105
use FILL  FILL_4593
timestamp 1711653199
transform 1 0 1024 0 1 370
box -8 -3 16 105
use FILL  FILL_4594
timestamp 1711653199
transform 1 0 1016 0 1 370
box -8 -3 16 105
use FILL  FILL_4595
timestamp 1711653199
transform 1 0 992 0 1 370
box -8 -3 16 105
use FILL  FILL_4596
timestamp 1711653199
transform 1 0 984 0 1 370
box -8 -3 16 105
use FILL  FILL_4597
timestamp 1711653199
transform 1 0 944 0 1 370
box -8 -3 16 105
use FILL  FILL_4598
timestamp 1711653199
transform 1 0 936 0 1 370
box -8 -3 16 105
use FILL  FILL_4599
timestamp 1711653199
transform 1 0 928 0 1 370
box -8 -3 16 105
use FILL  FILL_4600
timestamp 1711653199
transform 1 0 920 0 1 370
box -8 -3 16 105
use FILL  FILL_4601
timestamp 1711653199
transform 1 0 912 0 1 370
box -8 -3 16 105
use FILL  FILL_4602
timestamp 1711653199
transform 1 0 904 0 1 370
box -8 -3 16 105
use FILL  FILL_4603
timestamp 1711653199
transform 1 0 856 0 1 370
box -8 -3 16 105
use FILL  FILL_4604
timestamp 1711653199
transform 1 0 848 0 1 370
box -8 -3 16 105
use FILL  FILL_4605
timestamp 1711653199
transform 1 0 840 0 1 370
box -8 -3 16 105
use FILL  FILL_4606
timestamp 1711653199
transform 1 0 800 0 1 370
box -8 -3 16 105
use FILL  FILL_4607
timestamp 1711653199
transform 1 0 792 0 1 370
box -8 -3 16 105
use FILL  FILL_4608
timestamp 1711653199
transform 1 0 784 0 1 370
box -8 -3 16 105
use FILL  FILL_4609
timestamp 1711653199
transform 1 0 776 0 1 370
box -8 -3 16 105
use FILL  FILL_4610
timestamp 1711653199
transform 1 0 744 0 1 370
box -8 -3 16 105
use FILL  FILL_4611
timestamp 1711653199
transform 1 0 736 0 1 370
box -8 -3 16 105
use FILL  FILL_4612
timestamp 1711653199
transform 1 0 696 0 1 370
box -8 -3 16 105
use FILL  FILL_4613
timestamp 1711653199
transform 1 0 688 0 1 370
box -8 -3 16 105
use FILL  FILL_4614
timestamp 1711653199
transform 1 0 680 0 1 370
box -8 -3 16 105
use FILL  FILL_4615
timestamp 1711653199
transform 1 0 672 0 1 370
box -8 -3 16 105
use FILL  FILL_4616
timestamp 1711653199
transform 1 0 664 0 1 370
box -8 -3 16 105
use FILL  FILL_4617
timestamp 1711653199
transform 1 0 616 0 1 370
box -8 -3 16 105
use FILL  FILL_4618
timestamp 1711653199
transform 1 0 608 0 1 370
box -8 -3 16 105
use FILL  FILL_4619
timestamp 1711653199
transform 1 0 600 0 1 370
box -8 -3 16 105
use FILL  FILL_4620
timestamp 1711653199
transform 1 0 592 0 1 370
box -8 -3 16 105
use FILL  FILL_4621
timestamp 1711653199
transform 1 0 552 0 1 370
box -8 -3 16 105
use FILL  FILL_4622
timestamp 1711653199
transform 1 0 544 0 1 370
box -8 -3 16 105
use FILL  FILL_4623
timestamp 1711653199
transform 1 0 536 0 1 370
box -8 -3 16 105
use FILL  FILL_4624
timestamp 1711653199
transform 1 0 528 0 1 370
box -8 -3 16 105
use FILL  FILL_4625
timestamp 1711653199
transform 1 0 480 0 1 370
box -8 -3 16 105
use FILL  FILL_4626
timestamp 1711653199
transform 1 0 472 0 1 370
box -8 -3 16 105
use FILL  FILL_4627
timestamp 1711653199
transform 1 0 464 0 1 370
box -8 -3 16 105
use FILL  FILL_4628
timestamp 1711653199
transform 1 0 456 0 1 370
box -8 -3 16 105
use FILL  FILL_4629
timestamp 1711653199
transform 1 0 432 0 1 370
box -8 -3 16 105
use FILL  FILL_4630
timestamp 1711653199
transform 1 0 424 0 1 370
box -8 -3 16 105
use FILL  FILL_4631
timestamp 1711653199
transform 1 0 384 0 1 370
box -8 -3 16 105
use FILL  FILL_4632
timestamp 1711653199
transform 1 0 352 0 1 370
box -8 -3 16 105
use FILL  FILL_4633
timestamp 1711653199
transform 1 0 344 0 1 370
box -8 -3 16 105
use FILL  FILL_4634
timestamp 1711653199
transform 1 0 336 0 1 370
box -8 -3 16 105
use FILL  FILL_4635
timestamp 1711653199
transform 1 0 328 0 1 370
box -8 -3 16 105
use FILL  FILL_4636
timestamp 1711653199
transform 1 0 296 0 1 370
box -8 -3 16 105
use FILL  FILL_4637
timestamp 1711653199
transform 1 0 272 0 1 370
box -8 -3 16 105
use FILL  FILL_4638
timestamp 1711653199
transform 1 0 264 0 1 370
box -8 -3 16 105
use FILL  FILL_4639
timestamp 1711653199
transform 1 0 256 0 1 370
box -8 -3 16 105
use FILL  FILL_4640
timestamp 1711653199
transform 1 0 232 0 1 370
box -8 -3 16 105
use FILL  FILL_4641
timestamp 1711653199
transform 1 0 224 0 1 370
box -8 -3 16 105
use FILL  FILL_4642
timestamp 1711653199
transform 1 0 216 0 1 370
box -8 -3 16 105
use FILL  FILL_4643
timestamp 1711653199
transform 1 0 168 0 1 370
box -8 -3 16 105
use FILL  FILL_4644
timestamp 1711653199
transform 1 0 160 0 1 370
box -8 -3 16 105
use FILL  FILL_4645
timestamp 1711653199
transform 1 0 152 0 1 370
box -8 -3 16 105
use FILL  FILL_4646
timestamp 1711653199
transform 1 0 144 0 1 370
box -8 -3 16 105
use FILL  FILL_4647
timestamp 1711653199
transform 1 0 136 0 1 370
box -8 -3 16 105
use FILL  FILL_4648
timestamp 1711653199
transform 1 0 128 0 1 370
box -8 -3 16 105
use FILL  FILL_4649
timestamp 1711653199
transform 1 0 80 0 1 370
box -8 -3 16 105
use FILL  FILL_4650
timestamp 1711653199
transform 1 0 72 0 1 370
box -8 -3 16 105
use FILL  FILL_4651
timestamp 1711653199
transform 1 0 3392 0 -1 370
box -8 -3 16 105
use FILL  FILL_4652
timestamp 1711653199
transform 1 0 3384 0 -1 370
box -8 -3 16 105
use FILL  FILL_4653
timestamp 1711653199
transform 1 0 3344 0 -1 370
box -8 -3 16 105
use FILL  FILL_4654
timestamp 1711653199
transform 1 0 3336 0 -1 370
box -8 -3 16 105
use FILL  FILL_4655
timestamp 1711653199
transform 1 0 3328 0 -1 370
box -8 -3 16 105
use FILL  FILL_4656
timestamp 1711653199
transform 1 0 3320 0 -1 370
box -8 -3 16 105
use FILL  FILL_4657
timestamp 1711653199
transform 1 0 3272 0 -1 370
box -8 -3 16 105
use FILL  FILL_4658
timestamp 1711653199
transform 1 0 3264 0 -1 370
box -8 -3 16 105
use FILL  FILL_4659
timestamp 1711653199
transform 1 0 3256 0 -1 370
box -8 -3 16 105
use FILL  FILL_4660
timestamp 1711653199
transform 1 0 3248 0 -1 370
box -8 -3 16 105
use FILL  FILL_4661
timestamp 1711653199
transform 1 0 3240 0 -1 370
box -8 -3 16 105
use FILL  FILL_4662
timestamp 1711653199
transform 1 0 3232 0 -1 370
box -8 -3 16 105
use FILL  FILL_4663
timestamp 1711653199
transform 1 0 3200 0 -1 370
box -8 -3 16 105
use FILL  FILL_4664
timestamp 1711653199
transform 1 0 3192 0 -1 370
box -8 -3 16 105
use FILL  FILL_4665
timestamp 1711653199
transform 1 0 3184 0 -1 370
box -8 -3 16 105
use FILL  FILL_4666
timestamp 1711653199
transform 1 0 3144 0 -1 370
box -8 -3 16 105
use FILL  FILL_4667
timestamp 1711653199
transform 1 0 3136 0 -1 370
box -8 -3 16 105
use FILL  FILL_4668
timestamp 1711653199
transform 1 0 3128 0 -1 370
box -8 -3 16 105
use FILL  FILL_4669
timestamp 1711653199
transform 1 0 3120 0 -1 370
box -8 -3 16 105
use FILL  FILL_4670
timestamp 1711653199
transform 1 0 3112 0 -1 370
box -8 -3 16 105
use FILL  FILL_4671
timestamp 1711653199
transform 1 0 3104 0 -1 370
box -8 -3 16 105
use FILL  FILL_4672
timestamp 1711653199
transform 1 0 3080 0 -1 370
box -8 -3 16 105
use FILL  FILL_4673
timestamp 1711653199
transform 1 0 3072 0 -1 370
box -8 -3 16 105
use FILL  FILL_4674
timestamp 1711653199
transform 1 0 3032 0 -1 370
box -8 -3 16 105
use FILL  FILL_4675
timestamp 1711653199
transform 1 0 3024 0 -1 370
box -8 -3 16 105
use FILL  FILL_4676
timestamp 1711653199
transform 1 0 3016 0 -1 370
box -8 -3 16 105
use FILL  FILL_4677
timestamp 1711653199
transform 1 0 3008 0 -1 370
box -8 -3 16 105
use FILL  FILL_4678
timestamp 1711653199
transform 1 0 3000 0 -1 370
box -8 -3 16 105
use FILL  FILL_4679
timestamp 1711653199
transform 1 0 2992 0 -1 370
box -8 -3 16 105
use FILL  FILL_4680
timestamp 1711653199
transform 1 0 2936 0 -1 370
box -8 -3 16 105
use FILL  FILL_4681
timestamp 1711653199
transform 1 0 2928 0 -1 370
box -8 -3 16 105
use FILL  FILL_4682
timestamp 1711653199
transform 1 0 2920 0 -1 370
box -8 -3 16 105
use FILL  FILL_4683
timestamp 1711653199
transform 1 0 2912 0 -1 370
box -8 -3 16 105
use FILL  FILL_4684
timestamp 1711653199
transform 1 0 2904 0 -1 370
box -8 -3 16 105
use FILL  FILL_4685
timestamp 1711653199
transform 1 0 2896 0 -1 370
box -8 -3 16 105
use FILL  FILL_4686
timestamp 1711653199
transform 1 0 2824 0 -1 370
box -8 -3 16 105
use FILL  FILL_4687
timestamp 1711653199
transform 1 0 2816 0 -1 370
box -8 -3 16 105
use FILL  FILL_4688
timestamp 1711653199
transform 1 0 2808 0 -1 370
box -8 -3 16 105
use FILL  FILL_4689
timestamp 1711653199
transform 1 0 2800 0 -1 370
box -8 -3 16 105
use FILL  FILL_4690
timestamp 1711653199
transform 1 0 2792 0 -1 370
box -8 -3 16 105
use FILL  FILL_4691
timestamp 1711653199
transform 1 0 2784 0 -1 370
box -8 -3 16 105
use FILL  FILL_4692
timestamp 1711653199
transform 1 0 2728 0 -1 370
box -8 -3 16 105
use FILL  FILL_4693
timestamp 1711653199
transform 1 0 2720 0 -1 370
box -8 -3 16 105
use FILL  FILL_4694
timestamp 1711653199
transform 1 0 2712 0 -1 370
box -8 -3 16 105
use FILL  FILL_4695
timestamp 1711653199
transform 1 0 2688 0 -1 370
box -8 -3 16 105
use FILL  FILL_4696
timestamp 1711653199
transform 1 0 2680 0 -1 370
box -8 -3 16 105
use FILL  FILL_4697
timestamp 1711653199
transform 1 0 2672 0 -1 370
box -8 -3 16 105
use FILL  FILL_4698
timestamp 1711653199
transform 1 0 2616 0 -1 370
box -8 -3 16 105
use FILL  FILL_4699
timestamp 1711653199
transform 1 0 2608 0 -1 370
box -8 -3 16 105
use FILL  FILL_4700
timestamp 1711653199
transform 1 0 2600 0 -1 370
box -8 -3 16 105
use FILL  FILL_4701
timestamp 1711653199
transform 1 0 2592 0 -1 370
box -8 -3 16 105
use FILL  FILL_4702
timestamp 1711653199
transform 1 0 2584 0 -1 370
box -8 -3 16 105
use FILL  FILL_4703
timestamp 1711653199
transform 1 0 2576 0 -1 370
box -8 -3 16 105
use FILL  FILL_4704
timestamp 1711653199
transform 1 0 2528 0 -1 370
box -8 -3 16 105
use FILL  FILL_4705
timestamp 1711653199
transform 1 0 2520 0 -1 370
box -8 -3 16 105
use FILL  FILL_4706
timestamp 1711653199
transform 1 0 2512 0 -1 370
box -8 -3 16 105
use FILL  FILL_4707
timestamp 1711653199
transform 1 0 2504 0 -1 370
box -8 -3 16 105
use FILL  FILL_4708
timestamp 1711653199
transform 1 0 2456 0 -1 370
box -8 -3 16 105
use FILL  FILL_4709
timestamp 1711653199
transform 1 0 2448 0 -1 370
box -8 -3 16 105
use FILL  FILL_4710
timestamp 1711653199
transform 1 0 2440 0 -1 370
box -8 -3 16 105
use FILL  FILL_4711
timestamp 1711653199
transform 1 0 2432 0 -1 370
box -8 -3 16 105
use FILL  FILL_4712
timestamp 1711653199
transform 1 0 2424 0 -1 370
box -8 -3 16 105
use FILL  FILL_4713
timestamp 1711653199
transform 1 0 2384 0 -1 370
box -8 -3 16 105
use FILL  FILL_4714
timestamp 1711653199
transform 1 0 2376 0 -1 370
box -8 -3 16 105
use FILL  FILL_4715
timestamp 1711653199
transform 1 0 2368 0 -1 370
box -8 -3 16 105
use FILL  FILL_4716
timestamp 1711653199
transform 1 0 2360 0 -1 370
box -8 -3 16 105
use FILL  FILL_4717
timestamp 1711653199
transform 1 0 2352 0 -1 370
box -8 -3 16 105
use FILL  FILL_4718
timestamp 1711653199
transform 1 0 2312 0 -1 370
box -8 -3 16 105
use FILL  FILL_4719
timestamp 1711653199
transform 1 0 2304 0 -1 370
box -8 -3 16 105
use FILL  FILL_4720
timestamp 1711653199
transform 1 0 2296 0 -1 370
box -8 -3 16 105
use FILL  FILL_4721
timestamp 1711653199
transform 1 0 2288 0 -1 370
box -8 -3 16 105
use FILL  FILL_4722
timestamp 1711653199
transform 1 0 2248 0 -1 370
box -8 -3 16 105
use FILL  FILL_4723
timestamp 1711653199
transform 1 0 2240 0 -1 370
box -8 -3 16 105
use FILL  FILL_4724
timestamp 1711653199
transform 1 0 2232 0 -1 370
box -8 -3 16 105
use FILL  FILL_4725
timestamp 1711653199
transform 1 0 2224 0 -1 370
box -8 -3 16 105
use FILL  FILL_4726
timestamp 1711653199
transform 1 0 2216 0 -1 370
box -8 -3 16 105
use FILL  FILL_4727
timestamp 1711653199
transform 1 0 2192 0 -1 370
box -8 -3 16 105
use FILL  FILL_4728
timestamp 1711653199
transform 1 0 2184 0 -1 370
box -8 -3 16 105
use FILL  FILL_4729
timestamp 1711653199
transform 1 0 2144 0 -1 370
box -8 -3 16 105
use FILL  FILL_4730
timestamp 1711653199
transform 1 0 2136 0 -1 370
box -8 -3 16 105
use FILL  FILL_4731
timestamp 1711653199
transform 1 0 2128 0 -1 370
box -8 -3 16 105
use FILL  FILL_4732
timestamp 1711653199
transform 1 0 2120 0 -1 370
box -8 -3 16 105
use FILL  FILL_4733
timestamp 1711653199
transform 1 0 2112 0 -1 370
box -8 -3 16 105
use FILL  FILL_4734
timestamp 1711653199
transform 1 0 2104 0 -1 370
box -8 -3 16 105
use FILL  FILL_4735
timestamp 1711653199
transform 1 0 2064 0 -1 370
box -8 -3 16 105
use FILL  FILL_4736
timestamp 1711653199
transform 1 0 2056 0 -1 370
box -8 -3 16 105
use FILL  FILL_4737
timestamp 1711653199
transform 1 0 2048 0 -1 370
box -8 -3 16 105
use FILL  FILL_4738
timestamp 1711653199
transform 1 0 2040 0 -1 370
box -8 -3 16 105
use FILL  FILL_4739
timestamp 1711653199
transform 1 0 1992 0 -1 370
box -8 -3 16 105
use FILL  FILL_4740
timestamp 1711653199
transform 1 0 1984 0 -1 370
box -8 -3 16 105
use FILL  FILL_4741
timestamp 1711653199
transform 1 0 1976 0 -1 370
box -8 -3 16 105
use FILL  FILL_4742
timestamp 1711653199
transform 1 0 1968 0 -1 370
box -8 -3 16 105
use FILL  FILL_4743
timestamp 1711653199
transform 1 0 1960 0 -1 370
box -8 -3 16 105
use FILL  FILL_4744
timestamp 1711653199
transform 1 0 1952 0 -1 370
box -8 -3 16 105
use FILL  FILL_4745
timestamp 1711653199
transform 1 0 1928 0 -1 370
box -8 -3 16 105
use FILL  FILL_4746
timestamp 1711653199
transform 1 0 1888 0 -1 370
box -8 -3 16 105
use FILL  FILL_4747
timestamp 1711653199
transform 1 0 1880 0 -1 370
box -8 -3 16 105
use FILL  FILL_4748
timestamp 1711653199
transform 1 0 1872 0 -1 370
box -8 -3 16 105
use FILL  FILL_4749
timestamp 1711653199
transform 1 0 1864 0 -1 370
box -8 -3 16 105
use FILL  FILL_4750
timestamp 1711653199
transform 1 0 1856 0 -1 370
box -8 -3 16 105
use FILL  FILL_4751
timestamp 1711653199
transform 1 0 1848 0 -1 370
box -8 -3 16 105
use FILL  FILL_4752
timestamp 1711653199
transform 1 0 1840 0 -1 370
box -8 -3 16 105
use FILL  FILL_4753
timestamp 1711653199
transform 1 0 1792 0 -1 370
box -8 -3 16 105
use FILL  FILL_4754
timestamp 1711653199
transform 1 0 1784 0 -1 370
box -8 -3 16 105
use FILL  FILL_4755
timestamp 1711653199
transform 1 0 1776 0 -1 370
box -8 -3 16 105
use FILL  FILL_4756
timestamp 1711653199
transform 1 0 1768 0 -1 370
box -8 -3 16 105
use FILL  FILL_4757
timestamp 1711653199
transform 1 0 1736 0 -1 370
box -8 -3 16 105
use FILL  FILL_4758
timestamp 1711653199
transform 1 0 1728 0 -1 370
box -8 -3 16 105
use FILL  FILL_4759
timestamp 1711653199
transform 1 0 1720 0 -1 370
box -8 -3 16 105
use FILL  FILL_4760
timestamp 1711653199
transform 1 0 1712 0 -1 370
box -8 -3 16 105
use FILL  FILL_4761
timestamp 1711653199
transform 1 0 1704 0 -1 370
box -8 -3 16 105
use FILL  FILL_4762
timestamp 1711653199
transform 1 0 1696 0 -1 370
box -8 -3 16 105
use FILL  FILL_4763
timestamp 1711653199
transform 1 0 1688 0 -1 370
box -8 -3 16 105
use FILL  FILL_4764
timestamp 1711653199
transform 1 0 1640 0 -1 370
box -8 -3 16 105
use FILL  FILL_4765
timestamp 1711653199
transform 1 0 1632 0 -1 370
box -8 -3 16 105
use FILL  FILL_4766
timestamp 1711653199
transform 1 0 1624 0 -1 370
box -8 -3 16 105
use FILL  FILL_4767
timestamp 1711653199
transform 1 0 1616 0 -1 370
box -8 -3 16 105
use FILL  FILL_4768
timestamp 1711653199
transform 1 0 1608 0 -1 370
box -8 -3 16 105
use FILL  FILL_4769
timestamp 1711653199
transform 1 0 1600 0 -1 370
box -8 -3 16 105
use FILL  FILL_4770
timestamp 1711653199
transform 1 0 1560 0 -1 370
box -8 -3 16 105
use FILL  FILL_4771
timestamp 1711653199
transform 1 0 1552 0 -1 370
box -8 -3 16 105
use FILL  FILL_4772
timestamp 1711653199
transform 1 0 1544 0 -1 370
box -8 -3 16 105
use FILL  FILL_4773
timestamp 1711653199
transform 1 0 1512 0 -1 370
box -8 -3 16 105
use FILL  FILL_4774
timestamp 1711653199
transform 1 0 1504 0 -1 370
box -8 -3 16 105
use FILL  FILL_4775
timestamp 1711653199
transform 1 0 1496 0 -1 370
box -8 -3 16 105
use FILL  FILL_4776
timestamp 1711653199
transform 1 0 1488 0 -1 370
box -8 -3 16 105
use FILL  FILL_4777
timestamp 1711653199
transform 1 0 1480 0 -1 370
box -8 -3 16 105
use FILL  FILL_4778
timestamp 1711653199
transform 1 0 1448 0 -1 370
box -8 -3 16 105
use FILL  FILL_4779
timestamp 1711653199
transform 1 0 1416 0 -1 370
box -8 -3 16 105
use FILL  FILL_4780
timestamp 1711653199
transform 1 0 1408 0 -1 370
box -8 -3 16 105
use FILL  FILL_4781
timestamp 1711653199
transform 1 0 1400 0 -1 370
box -8 -3 16 105
use FILL  FILL_4782
timestamp 1711653199
transform 1 0 1392 0 -1 370
box -8 -3 16 105
use FILL  FILL_4783
timestamp 1711653199
transform 1 0 1384 0 -1 370
box -8 -3 16 105
use FILL  FILL_4784
timestamp 1711653199
transform 1 0 1376 0 -1 370
box -8 -3 16 105
use FILL  FILL_4785
timestamp 1711653199
transform 1 0 1344 0 -1 370
box -8 -3 16 105
use FILL  FILL_4786
timestamp 1711653199
transform 1 0 1336 0 -1 370
box -8 -3 16 105
use FILL  FILL_4787
timestamp 1711653199
transform 1 0 1304 0 -1 370
box -8 -3 16 105
use FILL  FILL_4788
timestamp 1711653199
transform 1 0 1296 0 -1 370
box -8 -3 16 105
use FILL  FILL_4789
timestamp 1711653199
transform 1 0 1288 0 -1 370
box -8 -3 16 105
use FILL  FILL_4790
timestamp 1711653199
transform 1 0 1280 0 -1 370
box -8 -3 16 105
use FILL  FILL_4791
timestamp 1711653199
transform 1 0 1272 0 -1 370
box -8 -3 16 105
use FILL  FILL_4792
timestamp 1711653199
transform 1 0 1232 0 -1 370
box -8 -3 16 105
use FILL  FILL_4793
timestamp 1711653199
transform 1 0 1224 0 -1 370
box -8 -3 16 105
use FILL  FILL_4794
timestamp 1711653199
transform 1 0 1216 0 -1 370
box -8 -3 16 105
use FILL  FILL_4795
timestamp 1711653199
transform 1 0 1208 0 -1 370
box -8 -3 16 105
use FILL  FILL_4796
timestamp 1711653199
transform 1 0 1168 0 -1 370
box -8 -3 16 105
use FILL  FILL_4797
timestamp 1711653199
transform 1 0 1160 0 -1 370
box -8 -3 16 105
use FILL  FILL_4798
timestamp 1711653199
transform 1 0 1136 0 -1 370
box -8 -3 16 105
use FILL  FILL_4799
timestamp 1711653199
transform 1 0 1128 0 -1 370
box -8 -3 16 105
use FILL  FILL_4800
timestamp 1711653199
transform 1 0 1120 0 -1 370
box -8 -3 16 105
use FILL  FILL_4801
timestamp 1711653199
transform 1 0 1112 0 -1 370
box -8 -3 16 105
use FILL  FILL_4802
timestamp 1711653199
transform 1 0 1072 0 -1 370
box -8 -3 16 105
use FILL  FILL_4803
timestamp 1711653199
transform 1 0 1064 0 -1 370
box -8 -3 16 105
use FILL  FILL_4804
timestamp 1711653199
transform 1 0 1056 0 -1 370
box -8 -3 16 105
use FILL  FILL_4805
timestamp 1711653199
transform 1 0 1008 0 -1 370
box -8 -3 16 105
use FILL  FILL_4806
timestamp 1711653199
transform 1 0 1000 0 -1 370
box -8 -3 16 105
use FILL  FILL_4807
timestamp 1711653199
transform 1 0 992 0 -1 370
box -8 -3 16 105
use FILL  FILL_4808
timestamp 1711653199
transform 1 0 984 0 -1 370
box -8 -3 16 105
use FILL  FILL_4809
timestamp 1711653199
transform 1 0 976 0 -1 370
box -8 -3 16 105
use FILL  FILL_4810
timestamp 1711653199
transform 1 0 928 0 -1 370
box -8 -3 16 105
use FILL  FILL_4811
timestamp 1711653199
transform 1 0 920 0 -1 370
box -8 -3 16 105
use FILL  FILL_4812
timestamp 1711653199
transform 1 0 912 0 -1 370
box -8 -3 16 105
use FILL  FILL_4813
timestamp 1711653199
transform 1 0 904 0 -1 370
box -8 -3 16 105
use FILL  FILL_4814
timestamp 1711653199
transform 1 0 864 0 -1 370
box -8 -3 16 105
use FILL  FILL_4815
timestamp 1711653199
transform 1 0 856 0 -1 370
box -8 -3 16 105
use FILL  FILL_4816
timestamp 1711653199
transform 1 0 816 0 -1 370
box -8 -3 16 105
use FILL  FILL_4817
timestamp 1711653199
transform 1 0 808 0 -1 370
box -8 -3 16 105
use FILL  FILL_4818
timestamp 1711653199
transform 1 0 800 0 -1 370
box -8 -3 16 105
use FILL  FILL_4819
timestamp 1711653199
transform 1 0 792 0 -1 370
box -8 -3 16 105
use FILL  FILL_4820
timestamp 1711653199
transform 1 0 768 0 -1 370
box -8 -3 16 105
use FILL  FILL_4821
timestamp 1711653199
transform 1 0 728 0 -1 370
box -8 -3 16 105
use FILL  FILL_4822
timestamp 1711653199
transform 1 0 720 0 -1 370
box -8 -3 16 105
use FILL  FILL_4823
timestamp 1711653199
transform 1 0 712 0 -1 370
box -8 -3 16 105
use FILL  FILL_4824
timestamp 1711653199
transform 1 0 704 0 -1 370
box -8 -3 16 105
use FILL  FILL_4825
timestamp 1711653199
transform 1 0 664 0 -1 370
box -8 -3 16 105
use FILL  FILL_4826
timestamp 1711653199
transform 1 0 656 0 -1 370
box -8 -3 16 105
use FILL  FILL_4827
timestamp 1711653199
transform 1 0 608 0 -1 370
box -8 -3 16 105
use FILL  FILL_4828
timestamp 1711653199
transform 1 0 600 0 -1 370
box -8 -3 16 105
use FILL  FILL_4829
timestamp 1711653199
transform 1 0 592 0 -1 370
box -8 -3 16 105
use FILL  FILL_4830
timestamp 1711653199
transform 1 0 584 0 -1 370
box -8 -3 16 105
use FILL  FILL_4831
timestamp 1711653199
transform 1 0 576 0 -1 370
box -8 -3 16 105
use FILL  FILL_4832
timestamp 1711653199
transform 1 0 536 0 -1 370
box -8 -3 16 105
use FILL  FILL_4833
timestamp 1711653199
transform 1 0 528 0 -1 370
box -8 -3 16 105
use FILL  FILL_4834
timestamp 1711653199
transform 1 0 488 0 -1 370
box -8 -3 16 105
use FILL  FILL_4835
timestamp 1711653199
transform 1 0 480 0 -1 370
box -8 -3 16 105
use FILL  FILL_4836
timestamp 1711653199
transform 1 0 472 0 -1 370
box -8 -3 16 105
use FILL  FILL_4837
timestamp 1711653199
transform 1 0 464 0 -1 370
box -8 -3 16 105
use FILL  FILL_4838
timestamp 1711653199
transform 1 0 456 0 -1 370
box -8 -3 16 105
use FILL  FILL_4839
timestamp 1711653199
transform 1 0 384 0 -1 370
box -8 -3 16 105
use FILL  FILL_4840
timestamp 1711653199
transform 1 0 376 0 -1 370
box -8 -3 16 105
use FILL  FILL_4841
timestamp 1711653199
transform 1 0 368 0 -1 370
box -8 -3 16 105
use FILL  FILL_4842
timestamp 1711653199
transform 1 0 360 0 -1 370
box -8 -3 16 105
use FILL  FILL_4843
timestamp 1711653199
transform 1 0 352 0 -1 370
box -8 -3 16 105
use FILL  FILL_4844
timestamp 1711653199
transform 1 0 344 0 -1 370
box -8 -3 16 105
use FILL  FILL_4845
timestamp 1711653199
transform 1 0 280 0 -1 370
box -8 -3 16 105
use FILL  FILL_4846
timestamp 1711653199
transform 1 0 272 0 -1 370
box -8 -3 16 105
use FILL  FILL_4847
timestamp 1711653199
transform 1 0 264 0 -1 370
box -8 -3 16 105
use FILL  FILL_4848
timestamp 1711653199
transform 1 0 224 0 -1 370
box -8 -3 16 105
use FILL  FILL_4849
timestamp 1711653199
transform 1 0 216 0 -1 370
box -8 -3 16 105
use FILL  FILL_4850
timestamp 1711653199
transform 1 0 184 0 -1 370
box -8 -3 16 105
use FILL  FILL_4851
timestamp 1711653199
transform 1 0 176 0 -1 370
box -8 -3 16 105
use FILL  FILL_4852
timestamp 1711653199
transform 1 0 168 0 -1 370
box -8 -3 16 105
use FILL  FILL_4853
timestamp 1711653199
transform 1 0 160 0 -1 370
box -8 -3 16 105
use FILL  FILL_4854
timestamp 1711653199
transform 1 0 128 0 -1 370
box -8 -3 16 105
use FILL  FILL_4855
timestamp 1711653199
transform 1 0 88 0 -1 370
box -8 -3 16 105
use FILL  FILL_4856
timestamp 1711653199
transform 1 0 80 0 -1 370
box -8 -3 16 105
use FILL  FILL_4857
timestamp 1711653199
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_4858
timestamp 1711653199
transform 1 0 3392 0 1 170
box -8 -3 16 105
use FILL  FILL_4859
timestamp 1711653199
transform 1 0 3384 0 1 170
box -8 -3 16 105
use FILL  FILL_4860
timestamp 1711653199
transform 1 0 3376 0 1 170
box -8 -3 16 105
use FILL  FILL_4861
timestamp 1711653199
transform 1 0 3368 0 1 170
box -8 -3 16 105
use FILL  FILL_4862
timestamp 1711653199
transform 1 0 3360 0 1 170
box -8 -3 16 105
use FILL  FILL_4863
timestamp 1711653199
transform 1 0 3352 0 1 170
box -8 -3 16 105
use FILL  FILL_4864
timestamp 1711653199
transform 1 0 3344 0 1 170
box -8 -3 16 105
use FILL  FILL_4865
timestamp 1711653199
transform 1 0 3336 0 1 170
box -8 -3 16 105
use FILL  FILL_4866
timestamp 1711653199
transform 1 0 3288 0 1 170
box -8 -3 16 105
use FILL  FILL_4867
timestamp 1711653199
transform 1 0 3280 0 1 170
box -8 -3 16 105
use FILL  FILL_4868
timestamp 1711653199
transform 1 0 3272 0 1 170
box -8 -3 16 105
use FILL  FILL_4869
timestamp 1711653199
transform 1 0 3240 0 1 170
box -8 -3 16 105
use FILL  FILL_4870
timestamp 1711653199
transform 1 0 3232 0 1 170
box -8 -3 16 105
use FILL  FILL_4871
timestamp 1711653199
transform 1 0 3224 0 1 170
box -8 -3 16 105
use FILL  FILL_4872
timestamp 1711653199
transform 1 0 3216 0 1 170
box -8 -3 16 105
use FILL  FILL_4873
timestamp 1711653199
transform 1 0 3208 0 1 170
box -8 -3 16 105
use FILL  FILL_4874
timestamp 1711653199
transform 1 0 3160 0 1 170
box -8 -3 16 105
use FILL  FILL_4875
timestamp 1711653199
transform 1 0 3152 0 1 170
box -8 -3 16 105
use FILL  FILL_4876
timestamp 1711653199
transform 1 0 3144 0 1 170
box -8 -3 16 105
use FILL  FILL_4877
timestamp 1711653199
transform 1 0 3136 0 1 170
box -8 -3 16 105
use FILL  FILL_4878
timestamp 1711653199
transform 1 0 3128 0 1 170
box -8 -3 16 105
use FILL  FILL_4879
timestamp 1711653199
transform 1 0 3080 0 1 170
box -8 -3 16 105
use FILL  FILL_4880
timestamp 1711653199
transform 1 0 3072 0 1 170
box -8 -3 16 105
use FILL  FILL_4881
timestamp 1711653199
transform 1 0 3064 0 1 170
box -8 -3 16 105
use FILL  FILL_4882
timestamp 1711653199
transform 1 0 3056 0 1 170
box -8 -3 16 105
use FILL  FILL_4883
timestamp 1711653199
transform 1 0 3024 0 1 170
box -8 -3 16 105
use FILL  FILL_4884
timestamp 1711653199
transform 1 0 3016 0 1 170
box -8 -3 16 105
use FILL  FILL_4885
timestamp 1711653199
transform 1 0 3008 0 1 170
box -8 -3 16 105
use FILL  FILL_4886
timestamp 1711653199
transform 1 0 3000 0 1 170
box -8 -3 16 105
use FILL  FILL_4887
timestamp 1711653199
transform 1 0 2952 0 1 170
box -8 -3 16 105
use FILL  FILL_4888
timestamp 1711653199
transform 1 0 2944 0 1 170
box -8 -3 16 105
use FILL  FILL_4889
timestamp 1711653199
transform 1 0 2936 0 1 170
box -8 -3 16 105
use FILL  FILL_4890
timestamp 1711653199
transform 1 0 2928 0 1 170
box -8 -3 16 105
use FILL  FILL_4891
timestamp 1711653199
transform 1 0 2888 0 1 170
box -8 -3 16 105
use FILL  FILL_4892
timestamp 1711653199
transform 1 0 2880 0 1 170
box -8 -3 16 105
use FILL  FILL_4893
timestamp 1711653199
transform 1 0 2872 0 1 170
box -8 -3 16 105
use FILL  FILL_4894
timestamp 1711653199
transform 1 0 2864 0 1 170
box -8 -3 16 105
use FILL  FILL_4895
timestamp 1711653199
transform 1 0 2840 0 1 170
box -8 -3 16 105
use FILL  FILL_4896
timestamp 1711653199
transform 1 0 2792 0 1 170
box -8 -3 16 105
use FILL  FILL_4897
timestamp 1711653199
transform 1 0 2784 0 1 170
box -8 -3 16 105
use FILL  FILL_4898
timestamp 1711653199
transform 1 0 2776 0 1 170
box -8 -3 16 105
use FILL  FILL_4899
timestamp 1711653199
transform 1 0 2768 0 1 170
box -8 -3 16 105
use FILL  FILL_4900
timestamp 1711653199
transform 1 0 2696 0 1 170
box -8 -3 16 105
use FILL  FILL_4901
timestamp 1711653199
transform 1 0 2688 0 1 170
box -8 -3 16 105
use FILL  FILL_4902
timestamp 1711653199
transform 1 0 2680 0 1 170
box -8 -3 16 105
use FILL  FILL_4903
timestamp 1711653199
transform 1 0 2672 0 1 170
box -8 -3 16 105
use FILL  FILL_4904
timestamp 1711653199
transform 1 0 2664 0 1 170
box -8 -3 16 105
use FILL  FILL_4905
timestamp 1711653199
transform 1 0 2624 0 1 170
box -8 -3 16 105
use FILL  FILL_4906
timestamp 1711653199
transform 1 0 2616 0 1 170
box -8 -3 16 105
use FILL  FILL_4907
timestamp 1711653199
transform 1 0 2608 0 1 170
box -8 -3 16 105
use FILL  FILL_4908
timestamp 1711653199
transform 1 0 2584 0 1 170
box -8 -3 16 105
use FILL  FILL_4909
timestamp 1711653199
transform 1 0 2576 0 1 170
box -8 -3 16 105
use FILL  FILL_4910
timestamp 1711653199
transform 1 0 2568 0 1 170
box -8 -3 16 105
use FILL  FILL_4911
timestamp 1711653199
transform 1 0 2560 0 1 170
box -8 -3 16 105
use FILL  FILL_4912
timestamp 1711653199
transform 1 0 2520 0 1 170
box -8 -3 16 105
use FILL  FILL_4913
timestamp 1711653199
transform 1 0 2512 0 1 170
box -8 -3 16 105
use FILL  FILL_4914
timestamp 1711653199
transform 1 0 2504 0 1 170
box -8 -3 16 105
use FILL  FILL_4915
timestamp 1711653199
transform 1 0 2496 0 1 170
box -8 -3 16 105
use FILL  FILL_4916
timestamp 1711653199
transform 1 0 2488 0 1 170
box -8 -3 16 105
use FILL  FILL_4917
timestamp 1711653199
transform 1 0 2480 0 1 170
box -8 -3 16 105
use FILL  FILL_4918
timestamp 1711653199
transform 1 0 2432 0 1 170
box -8 -3 16 105
use FILL  FILL_4919
timestamp 1711653199
transform 1 0 2424 0 1 170
box -8 -3 16 105
use FILL  FILL_4920
timestamp 1711653199
transform 1 0 2416 0 1 170
box -8 -3 16 105
use FILL  FILL_4921
timestamp 1711653199
transform 1 0 2408 0 1 170
box -8 -3 16 105
use FILL  FILL_4922
timestamp 1711653199
transform 1 0 2400 0 1 170
box -8 -3 16 105
use FILL  FILL_4923
timestamp 1711653199
transform 1 0 2360 0 1 170
box -8 -3 16 105
use FILL  FILL_4924
timestamp 1711653199
transform 1 0 2352 0 1 170
box -8 -3 16 105
use FILL  FILL_4925
timestamp 1711653199
transform 1 0 2344 0 1 170
box -8 -3 16 105
use FILL  FILL_4926
timestamp 1711653199
transform 1 0 2336 0 1 170
box -8 -3 16 105
use FILL  FILL_4927
timestamp 1711653199
transform 1 0 2296 0 1 170
box -8 -3 16 105
use FILL  FILL_4928
timestamp 1711653199
transform 1 0 2288 0 1 170
box -8 -3 16 105
use FILL  FILL_4929
timestamp 1711653199
transform 1 0 2280 0 1 170
box -8 -3 16 105
use FILL  FILL_4930
timestamp 1711653199
transform 1 0 2272 0 1 170
box -8 -3 16 105
use FILL  FILL_4931
timestamp 1711653199
transform 1 0 2264 0 1 170
box -8 -3 16 105
use FILL  FILL_4932
timestamp 1711653199
transform 1 0 2224 0 1 170
box -8 -3 16 105
use FILL  FILL_4933
timestamp 1711653199
transform 1 0 2216 0 1 170
box -8 -3 16 105
use FILL  FILL_4934
timestamp 1711653199
transform 1 0 2208 0 1 170
box -8 -3 16 105
use FILL  FILL_4935
timestamp 1711653199
transform 1 0 2200 0 1 170
box -8 -3 16 105
use FILL  FILL_4936
timestamp 1711653199
transform 1 0 2192 0 1 170
box -8 -3 16 105
use FILL  FILL_4937
timestamp 1711653199
transform 1 0 2152 0 1 170
box -8 -3 16 105
use FILL  FILL_4938
timestamp 1711653199
transform 1 0 2144 0 1 170
box -8 -3 16 105
use FILL  FILL_4939
timestamp 1711653199
transform 1 0 2136 0 1 170
box -8 -3 16 105
use FILL  FILL_4940
timestamp 1711653199
transform 1 0 2128 0 1 170
box -8 -3 16 105
use FILL  FILL_4941
timestamp 1711653199
transform 1 0 2120 0 1 170
box -8 -3 16 105
use FILL  FILL_4942
timestamp 1711653199
transform 1 0 2080 0 1 170
box -8 -3 16 105
use FILL  FILL_4943
timestamp 1711653199
transform 1 0 2072 0 1 170
box -8 -3 16 105
use FILL  FILL_4944
timestamp 1711653199
transform 1 0 2064 0 1 170
box -8 -3 16 105
use FILL  FILL_4945
timestamp 1711653199
transform 1 0 2056 0 1 170
box -8 -3 16 105
use FILL  FILL_4946
timestamp 1711653199
transform 1 0 2048 0 1 170
box -8 -3 16 105
use FILL  FILL_4947
timestamp 1711653199
transform 1 0 2040 0 1 170
box -8 -3 16 105
use FILL  FILL_4948
timestamp 1711653199
transform 1 0 2000 0 1 170
box -8 -3 16 105
use FILL  FILL_4949
timestamp 1711653199
transform 1 0 1992 0 1 170
box -8 -3 16 105
use FILL  FILL_4950
timestamp 1711653199
transform 1 0 1984 0 1 170
box -8 -3 16 105
use FILL  FILL_4951
timestamp 1711653199
transform 1 0 1976 0 1 170
box -8 -3 16 105
use FILL  FILL_4952
timestamp 1711653199
transform 1 0 1944 0 1 170
box -8 -3 16 105
use FILL  FILL_4953
timestamp 1711653199
transform 1 0 1936 0 1 170
box -8 -3 16 105
use FILL  FILL_4954
timestamp 1711653199
transform 1 0 1928 0 1 170
box -8 -3 16 105
use FILL  FILL_4955
timestamp 1711653199
transform 1 0 1920 0 1 170
box -8 -3 16 105
use FILL  FILL_4956
timestamp 1711653199
transform 1 0 1912 0 1 170
box -8 -3 16 105
use FILL  FILL_4957
timestamp 1711653199
transform 1 0 1880 0 1 170
box -8 -3 16 105
use FILL  FILL_4958
timestamp 1711653199
transform 1 0 1872 0 1 170
box -8 -3 16 105
use FILL  FILL_4959
timestamp 1711653199
transform 1 0 1864 0 1 170
box -8 -3 16 105
use FILL  FILL_4960
timestamp 1711653199
transform 1 0 1856 0 1 170
box -8 -3 16 105
use FILL  FILL_4961
timestamp 1711653199
transform 1 0 1824 0 1 170
box -8 -3 16 105
use FILL  FILL_4962
timestamp 1711653199
transform 1 0 1816 0 1 170
box -8 -3 16 105
use FILL  FILL_4963
timestamp 1711653199
transform 1 0 1808 0 1 170
box -8 -3 16 105
use FILL  FILL_4964
timestamp 1711653199
transform 1 0 1800 0 1 170
box -8 -3 16 105
use FILL  FILL_4965
timestamp 1711653199
transform 1 0 1792 0 1 170
box -8 -3 16 105
use FILL  FILL_4966
timestamp 1711653199
transform 1 0 1784 0 1 170
box -8 -3 16 105
use FILL  FILL_4967
timestamp 1711653199
transform 1 0 1752 0 1 170
box -8 -3 16 105
use FILL  FILL_4968
timestamp 1711653199
transform 1 0 1728 0 1 170
box -8 -3 16 105
use FILL  FILL_4969
timestamp 1711653199
transform 1 0 1720 0 1 170
box -8 -3 16 105
use FILL  FILL_4970
timestamp 1711653199
transform 1 0 1712 0 1 170
box -8 -3 16 105
use FILL  FILL_4971
timestamp 1711653199
transform 1 0 1704 0 1 170
box -8 -3 16 105
use FILL  FILL_4972
timestamp 1711653199
transform 1 0 1696 0 1 170
box -8 -3 16 105
use FILL  FILL_4973
timestamp 1711653199
transform 1 0 1688 0 1 170
box -8 -3 16 105
use FILL  FILL_4974
timestamp 1711653199
transform 1 0 1680 0 1 170
box -8 -3 16 105
use FILL  FILL_4975
timestamp 1711653199
transform 1 0 1672 0 1 170
box -8 -3 16 105
use FILL  FILL_4976
timestamp 1711653199
transform 1 0 1624 0 1 170
box -8 -3 16 105
use FILL  FILL_4977
timestamp 1711653199
transform 1 0 1616 0 1 170
box -8 -3 16 105
use FILL  FILL_4978
timestamp 1711653199
transform 1 0 1608 0 1 170
box -8 -3 16 105
use FILL  FILL_4979
timestamp 1711653199
transform 1 0 1600 0 1 170
box -8 -3 16 105
use FILL  FILL_4980
timestamp 1711653199
transform 1 0 1592 0 1 170
box -8 -3 16 105
use FILL  FILL_4981
timestamp 1711653199
transform 1 0 1584 0 1 170
box -8 -3 16 105
use FILL  FILL_4982
timestamp 1711653199
transform 1 0 1576 0 1 170
box -8 -3 16 105
use FILL  FILL_4983
timestamp 1711653199
transform 1 0 1568 0 1 170
box -8 -3 16 105
use FILL  FILL_4984
timestamp 1711653199
transform 1 0 1544 0 1 170
box -8 -3 16 105
use FILL  FILL_4985
timestamp 1711653199
transform 1 0 1536 0 1 170
box -8 -3 16 105
use FILL  FILL_4986
timestamp 1711653199
transform 1 0 1528 0 1 170
box -8 -3 16 105
use FILL  FILL_4987
timestamp 1711653199
transform 1 0 1520 0 1 170
box -8 -3 16 105
use FILL  FILL_4988
timestamp 1711653199
transform 1 0 1488 0 1 170
box -8 -3 16 105
use FILL  FILL_4989
timestamp 1711653199
transform 1 0 1480 0 1 170
box -8 -3 16 105
use FILL  FILL_4990
timestamp 1711653199
transform 1 0 1472 0 1 170
box -8 -3 16 105
use FILL  FILL_4991
timestamp 1711653199
transform 1 0 1464 0 1 170
box -8 -3 16 105
use FILL  FILL_4992
timestamp 1711653199
transform 1 0 1456 0 1 170
box -8 -3 16 105
use FILL  FILL_4993
timestamp 1711653199
transform 1 0 1448 0 1 170
box -8 -3 16 105
use FILL  FILL_4994
timestamp 1711653199
transform 1 0 1416 0 1 170
box -8 -3 16 105
use FILL  FILL_4995
timestamp 1711653199
transform 1 0 1408 0 1 170
box -8 -3 16 105
use FILL  FILL_4996
timestamp 1711653199
transform 1 0 1400 0 1 170
box -8 -3 16 105
use FILL  FILL_4997
timestamp 1711653199
transform 1 0 1392 0 1 170
box -8 -3 16 105
use FILL  FILL_4998
timestamp 1711653199
transform 1 0 1384 0 1 170
box -8 -3 16 105
use FILL  FILL_4999
timestamp 1711653199
transform 1 0 1376 0 1 170
box -8 -3 16 105
use FILL  FILL_5000
timestamp 1711653199
transform 1 0 1368 0 1 170
box -8 -3 16 105
use FILL  FILL_5001
timestamp 1711653199
transform 1 0 1320 0 1 170
box -8 -3 16 105
use FILL  FILL_5002
timestamp 1711653199
transform 1 0 1312 0 1 170
box -8 -3 16 105
use FILL  FILL_5003
timestamp 1711653199
transform 1 0 1304 0 1 170
box -8 -3 16 105
use FILL  FILL_5004
timestamp 1711653199
transform 1 0 1296 0 1 170
box -8 -3 16 105
use FILL  FILL_5005
timestamp 1711653199
transform 1 0 1288 0 1 170
box -8 -3 16 105
use FILL  FILL_5006
timestamp 1711653199
transform 1 0 1280 0 1 170
box -8 -3 16 105
use FILL  FILL_5007
timestamp 1711653199
transform 1 0 1272 0 1 170
box -8 -3 16 105
use FILL  FILL_5008
timestamp 1711653199
transform 1 0 1232 0 1 170
box -8 -3 16 105
use FILL  FILL_5009
timestamp 1711653199
transform 1 0 1224 0 1 170
box -8 -3 16 105
use FILL  FILL_5010
timestamp 1711653199
transform 1 0 1216 0 1 170
box -8 -3 16 105
use FILL  FILL_5011
timestamp 1711653199
transform 1 0 1208 0 1 170
box -8 -3 16 105
use FILL  FILL_5012
timestamp 1711653199
transform 1 0 1200 0 1 170
box -8 -3 16 105
use FILL  FILL_5013
timestamp 1711653199
transform 1 0 1192 0 1 170
box -8 -3 16 105
use FILL  FILL_5014
timestamp 1711653199
transform 1 0 1184 0 1 170
box -8 -3 16 105
use FILL  FILL_5015
timestamp 1711653199
transform 1 0 1144 0 1 170
box -8 -3 16 105
use FILL  FILL_5016
timestamp 1711653199
transform 1 0 1136 0 1 170
box -8 -3 16 105
use FILL  FILL_5017
timestamp 1711653199
transform 1 0 1128 0 1 170
box -8 -3 16 105
use FILL  FILL_5018
timestamp 1711653199
transform 1 0 1120 0 1 170
box -8 -3 16 105
use FILL  FILL_5019
timestamp 1711653199
transform 1 0 1112 0 1 170
box -8 -3 16 105
use FILL  FILL_5020
timestamp 1711653199
transform 1 0 1104 0 1 170
box -8 -3 16 105
use FILL  FILL_5021
timestamp 1711653199
transform 1 0 1080 0 1 170
box -8 -3 16 105
use FILL  FILL_5022
timestamp 1711653199
transform 1 0 1072 0 1 170
box -8 -3 16 105
use FILL  FILL_5023
timestamp 1711653199
transform 1 0 1064 0 1 170
box -8 -3 16 105
use FILL  FILL_5024
timestamp 1711653199
transform 1 0 1056 0 1 170
box -8 -3 16 105
use FILL  FILL_5025
timestamp 1711653199
transform 1 0 1016 0 1 170
box -8 -3 16 105
use FILL  FILL_5026
timestamp 1711653199
transform 1 0 1008 0 1 170
box -8 -3 16 105
use FILL  FILL_5027
timestamp 1711653199
transform 1 0 1000 0 1 170
box -8 -3 16 105
use FILL  FILL_5028
timestamp 1711653199
transform 1 0 992 0 1 170
box -8 -3 16 105
use FILL  FILL_5029
timestamp 1711653199
transform 1 0 984 0 1 170
box -8 -3 16 105
use FILL  FILL_5030
timestamp 1711653199
transform 1 0 976 0 1 170
box -8 -3 16 105
use FILL  FILL_5031
timestamp 1711653199
transform 1 0 968 0 1 170
box -8 -3 16 105
use FILL  FILL_5032
timestamp 1711653199
transform 1 0 936 0 1 170
box -8 -3 16 105
use FILL  FILL_5033
timestamp 1711653199
transform 1 0 928 0 1 170
box -8 -3 16 105
use FILL  FILL_5034
timestamp 1711653199
transform 1 0 920 0 1 170
box -8 -3 16 105
use FILL  FILL_5035
timestamp 1711653199
transform 1 0 912 0 1 170
box -8 -3 16 105
use FILL  FILL_5036
timestamp 1711653199
transform 1 0 904 0 1 170
box -8 -3 16 105
use FILL  FILL_5037
timestamp 1711653199
transform 1 0 896 0 1 170
box -8 -3 16 105
use FILL  FILL_5038
timestamp 1711653199
transform 1 0 848 0 1 170
box -8 -3 16 105
use FILL  FILL_5039
timestamp 1711653199
transform 1 0 840 0 1 170
box -8 -3 16 105
use FILL  FILL_5040
timestamp 1711653199
transform 1 0 832 0 1 170
box -8 -3 16 105
use FILL  FILL_5041
timestamp 1711653199
transform 1 0 824 0 1 170
box -8 -3 16 105
use FILL  FILL_5042
timestamp 1711653199
transform 1 0 816 0 1 170
box -8 -3 16 105
use FILL  FILL_5043
timestamp 1711653199
transform 1 0 784 0 1 170
box -8 -3 16 105
use FILL  FILL_5044
timestamp 1711653199
transform 1 0 776 0 1 170
box -8 -3 16 105
use FILL  FILL_5045
timestamp 1711653199
transform 1 0 768 0 1 170
box -8 -3 16 105
use FILL  FILL_5046
timestamp 1711653199
transform 1 0 760 0 1 170
box -8 -3 16 105
use FILL  FILL_5047
timestamp 1711653199
transform 1 0 752 0 1 170
box -8 -3 16 105
use FILL  FILL_5048
timestamp 1711653199
transform 1 0 744 0 1 170
box -8 -3 16 105
use FILL  FILL_5049
timestamp 1711653199
transform 1 0 704 0 1 170
box -8 -3 16 105
use FILL  FILL_5050
timestamp 1711653199
transform 1 0 696 0 1 170
box -8 -3 16 105
use FILL  FILL_5051
timestamp 1711653199
transform 1 0 688 0 1 170
box -8 -3 16 105
use FILL  FILL_5052
timestamp 1711653199
transform 1 0 664 0 1 170
box -8 -3 16 105
use FILL  FILL_5053
timestamp 1711653199
transform 1 0 656 0 1 170
box -8 -3 16 105
use FILL  FILL_5054
timestamp 1711653199
transform 1 0 648 0 1 170
box -8 -3 16 105
use FILL  FILL_5055
timestamp 1711653199
transform 1 0 640 0 1 170
box -8 -3 16 105
use FILL  FILL_5056
timestamp 1711653199
transform 1 0 592 0 1 170
box -8 -3 16 105
use FILL  FILL_5057
timestamp 1711653199
transform 1 0 584 0 1 170
box -8 -3 16 105
use FILL  FILL_5058
timestamp 1711653199
transform 1 0 576 0 1 170
box -8 -3 16 105
use FILL  FILL_5059
timestamp 1711653199
transform 1 0 568 0 1 170
box -8 -3 16 105
use FILL  FILL_5060
timestamp 1711653199
transform 1 0 560 0 1 170
box -8 -3 16 105
use FILL  FILL_5061
timestamp 1711653199
transform 1 0 552 0 1 170
box -8 -3 16 105
use FILL  FILL_5062
timestamp 1711653199
transform 1 0 520 0 1 170
box -8 -3 16 105
use FILL  FILL_5063
timestamp 1711653199
transform 1 0 512 0 1 170
box -8 -3 16 105
use FILL  FILL_5064
timestamp 1711653199
transform 1 0 504 0 1 170
box -8 -3 16 105
use FILL  FILL_5065
timestamp 1711653199
transform 1 0 464 0 1 170
box -8 -3 16 105
use FILL  FILL_5066
timestamp 1711653199
transform 1 0 456 0 1 170
box -8 -3 16 105
use FILL  FILL_5067
timestamp 1711653199
transform 1 0 448 0 1 170
box -8 -3 16 105
use FILL  FILL_5068
timestamp 1711653199
transform 1 0 440 0 1 170
box -8 -3 16 105
use FILL  FILL_5069
timestamp 1711653199
transform 1 0 432 0 1 170
box -8 -3 16 105
use FILL  FILL_5070
timestamp 1711653199
transform 1 0 400 0 1 170
box -8 -3 16 105
use FILL  FILL_5071
timestamp 1711653199
transform 1 0 392 0 1 170
box -8 -3 16 105
use FILL  FILL_5072
timestamp 1711653199
transform 1 0 384 0 1 170
box -8 -3 16 105
use FILL  FILL_5073
timestamp 1711653199
transform 1 0 376 0 1 170
box -8 -3 16 105
use FILL  FILL_5074
timestamp 1711653199
transform 1 0 328 0 1 170
box -8 -3 16 105
use FILL  FILL_5075
timestamp 1711653199
transform 1 0 320 0 1 170
box -8 -3 16 105
use FILL  FILL_5076
timestamp 1711653199
transform 1 0 312 0 1 170
box -8 -3 16 105
use FILL  FILL_5077
timestamp 1711653199
transform 1 0 304 0 1 170
box -8 -3 16 105
use FILL  FILL_5078
timestamp 1711653199
transform 1 0 296 0 1 170
box -8 -3 16 105
use FILL  FILL_5079
timestamp 1711653199
transform 1 0 288 0 1 170
box -8 -3 16 105
use FILL  FILL_5080
timestamp 1711653199
transform 1 0 280 0 1 170
box -8 -3 16 105
use FILL  FILL_5081
timestamp 1711653199
transform 1 0 240 0 1 170
box -8 -3 16 105
use FILL  FILL_5082
timestamp 1711653199
transform 1 0 232 0 1 170
box -8 -3 16 105
use FILL  FILL_5083
timestamp 1711653199
transform 1 0 224 0 1 170
box -8 -3 16 105
use FILL  FILL_5084
timestamp 1711653199
transform 1 0 216 0 1 170
box -8 -3 16 105
use FILL  FILL_5085
timestamp 1711653199
transform 1 0 176 0 1 170
box -8 -3 16 105
use FILL  FILL_5086
timestamp 1711653199
transform 1 0 168 0 1 170
box -8 -3 16 105
use FILL  FILL_5087
timestamp 1711653199
transform 1 0 160 0 1 170
box -8 -3 16 105
use FILL  FILL_5088
timestamp 1711653199
transform 1 0 152 0 1 170
box -8 -3 16 105
use FILL  FILL_5089
timestamp 1711653199
transform 1 0 144 0 1 170
box -8 -3 16 105
use FILL  FILL_5090
timestamp 1711653199
transform 1 0 136 0 1 170
box -8 -3 16 105
use FILL  FILL_5091
timestamp 1711653199
transform 1 0 88 0 1 170
box -8 -3 16 105
use FILL  FILL_5092
timestamp 1711653199
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_5093
timestamp 1711653199
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_5094
timestamp 1711653199
transform 1 0 3392 0 -1 170
box -8 -3 16 105
use FILL  FILL_5095
timestamp 1711653199
transform 1 0 3384 0 -1 170
box -8 -3 16 105
use FILL  FILL_5096
timestamp 1711653199
transform 1 0 3376 0 -1 170
box -8 -3 16 105
use FILL  FILL_5097
timestamp 1711653199
transform 1 0 3368 0 -1 170
box -8 -3 16 105
use FILL  FILL_5098
timestamp 1711653199
transform 1 0 3360 0 -1 170
box -8 -3 16 105
use FILL  FILL_5099
timestamp 1711653199
transform 1 0 3352 0 -1 170
box -8 -3 16 105
use FILL  FILL_5100
timestamp 1711653199
transform 1 0 3344 0 -1 170
box -8 -3 16 105
use FILL  FILL_5101
timestamp 1711653199
transform 1 0 3336 0 -1 170
box -8 -3 16 105
use FILL  FILL_5102
timestamp 1711653199
transform 1 0 3328 0 -1 170
box -8 -3 16 105
use FILL  FILL_5103
timestamp 1711653199
transform 1 0 3280 0 -1 170
box -8 -3 16 105
use FILL  FILL_5104
timestamp 1711653199
transform 1 0 3272 0 -1 170
box -8 -3 16 105
use FILL  FILL_5105
timestamp 1711653199
transform 1 0 3264 0 -1 170
box -8 -3 16 105
use FILL  FILL_5106
timestamp 1711653199
transform 1 0 3256 0 -1 170
box -8 -3 16 105
use FILL  FILL_5107
timestamp 1711653199
transform 1 0 3248 0 -1 170
box -8 -3 16 105
use FILL  FILL_5108
timestamp 1711653199
transform 1 0 3240 0 -1 170
box -8 -3 16 105
use FILL  FILL_5109
timestamp 1711653199
transform 1 0 3232 0 -1 170
box -8 -3 16 105
use FILL  FILL_5110
timestamp 1711653199
transform 1 0 3224 0 -1 170
box -8 -3 16 105
use FILL  FILL_5111
timestamp 1711653199
transform 1 0 3216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5112
timestamp 1711653199
transform 1 0 3208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5113
timestamp 1711653199
transform 1 0 3160 0 -1 170
box -8 -3 16 105
use FILL  FILL_5114
timestamp 1711653199
transform 1 0 3152 0 -1 170
box -8 -3 16 105
use FILL  FILL_5115
timestamp 1711653199
transform 1 0 3144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5116
timestamp 1711653199
transform 1 0 3136 0 -1 170
box -8 -3 16 105
use FILL  FILL_5117
timestamp 1711653199
transform 1 0 3128 0 -1 170
box -8 -3 16 105
use FILL  FILL_5118
timestamp 1711653199
transform 1 0 3120 0 -1 170
box -8 -3 16 105
use FILL  FILL_5119
timestamp 1711653199
transform 1 0 3112 0 -1 170
box -8 -3 16 105
use FILL  FILL_5120
timestamp 1711653199
transform 1 0 3104 0 -1 170
box -8 -3 16 105
use FILL  FILL_5121
timestamp 1711653199
transform 1 0 3048 0 -1 170
box -8 -3 16 105
use FILL  FILL_5122
timestamp 1711653199
transform 1 0 3040 0 -1 170
box -8 -3 16 105
use FILL  FILL_5123
timestamp 1711653199
transform 1 0 3032 0 -1 170
box -8 -3 16 105
use FILL  FILL_5124
timestamp 1711653199
transform 1 0 3024 0 -1 170
box -8 -3 16 105
use FILL  FILL_5125
timestamp 1711653199
transform 1 0 3016 0 -1 170
box -8 -3 16 105
use FILL  FILL_5126
timestamp 1711653199
transform 1 0 3008 0 -1 170
box -8 -3 16 105
use FILL  FILL_5127
timestamp 1711653199
transform 1 0 3000 0 -1 170
box -8 -3 16 105
use FILL  FILL_5128
timestamp 1711653199
transform 1 0 2992 0 -1 170
box -8 -3 16 105
use FILL  FILL_5129
timestamp 1711653199
transform 1 0 2936 0 -1 170
box -8 -3 16 105
use FILL  FILL_5130
timestamp 1711653199
transform 1 0 2928 0 -1 170
box -8 -3 16 105
use FILL  FILL_5131
timestamp 1711653199
transform 1 0 2920 0 -1 170
box -8 -3 16 105
use FILL  FILL_5132
timestamp 1711653199
transform 1 0 2912 0 -1 170
box -8 -3 16 105
use FILL  FILL_5133
timestamp 1711653199
transform 1 0 2904 0 -1 170
box -8 -3 16 105
use FILL  FILL_5134
timestamp 1711653199
transform 1 0 2896 0 -1 170
box -8 -3 16 105
use FILL  FILL_5135
timestamp 1711653199
transform 1 0 2888 0 -1 170
box -8 -3 16 105
use FILL  FILL_5136
timestamp 1711653199
transform 1 0 2880 0 -1 170
box -8 -3 16 105
use FILL  FILL_5137
timestamp 1711653199
transform 1 0 2832 0 -1 170
box -8 -3 16 105
use FILL  FILL_5138
timestamp 1711653199
transform 1 0 2824 0 -1 170
box -8 -3 16 105
use FILL  FILL_5139
timestamp 1711653199
transform 1 0 2816 0 -1 170
box -8 -3 16 105
use FILL  FILL_5140
timestamp 1711653199
transform 1 0 2792 0 -1 170
box -8 -3 16 105
use FILL  FILL_5141
timestamp 1711653199
transform 1 0 2784 0 -1 170
box -8 -3 16 105
use FILL  FILL_5142
timestamp 1711653199
transform 1 0 2776 0 -1 170
box -8 -3 16 105
use FILL  FILL_5143
timestamp 1711653199
transform 1 0 2768 0 -1 170
box -8 -3 16 105
use FILL  FILL_5144
timestamp 1711653199
transform 1 0 2736 0 -1 170
box -8 -3 16 105
use FILL  FILL_5145
timestamp 1711653199
transform 1 0 2712 0 -1 170
box -8 -3 16 105
use FILL  FILL_5146
timestamp 1711653199
transform 1 0 2704 0 -1 170
box -8 -3 16 105
use FILL  FILL_5147
timestamp 1711653199
transform 1 0 2696 0 -1 170
box -8 -3 16 105
use FILL  FILL_5148
timestamp 1711653199
transform 1 0 2688 0 -1 170
box -8 -3 16 105
use FILL  FILL_5149
timestamp 1711653199
transform 1 0 2680 0 -1 170
box -8 -3 16 105
use FILL  FILL_5150
timestamp 1711653199
transform 1 0 2648 0 -1 170
box -8 -3 16 105
use FILL  FILL_5151
timestamp 1711653199
transform 1 0 2640 0 -1 170
box -8 -3 16 105
use FILL  FILL_5152
timestamp 1711653199
transform 1 0 2632 0 -1 170
box -8 -3 16 105
use FILL  FILL_5153
timestamp 1711653199
transform 1 0 2624 0 -1 170
box -8 -3 16 105
use FILL  FILL_5154
timestamp 1711653199
transform 1 0 2584 0 -1 170
box -8 -3 16 105
use FILL  FILL_5155
timestamp 1711653199
transform 1 0 2576 0 -1 170
box -8 -3 16 105
use FILL  FILL_5156
timestamp 1711653199
transform 1 0 2568 0 -1 170
box -8 -3 16 105
use FILL  FILL_5157
timestamp 1711653199
transform 1 0 2560 0 -1 170
box -8 -3 16 105
use FILL  FILL_5158
timestamp 1711653199
transform 1 0 2552 0 -1 170
box -8 -3 16 105
use FILL  FILL_5159
timestamp 1711653199
transform 1 0 2512 0 -1 170
box -8 -3 16 105
use FILL  FILL_5160
timestamp 1711653199
transform 1 0 2504 0 -1 170
box -8 -3 16 105
use FILL  FILL_5161
timestamp 1711653199
transform 1 0 2496 0 -1 170
box -8 -3 16 105
use FILL  FILL_5162
timestamp 1711653199
transform 1 0 2472 0 -1 170
box -8 -3 16 105
use FILL  FILL_5163
timestamp 1711653199
transform 1 0 2464 0 -1 170
box -8 -3 16 105
use FILL  FILL_5164
timestamp 1711653199
transform 1 0 2456 0 -1 170
box -8 -3 16 105
use FILL  FILL_5165
timestamp 1711653199
transform 1 0 2432 0 -1 170
box -8 -3 16 105
use FILL  FILL_5166
timestamp 1711653199
transform 1 0 2424 0 -1 170
box -8 -3 16 105
use FILL  FILL_5167
timestamp 1711653199
transform 1 0 2416 0 -1 170
box -8 -3 16 105
use FILL  FILL_5168
timestamp 1711653199
transform 1 0 2408 0 -1 170
box -8 -3 16 105
use FILL  FILL_5169
timestamp 1711653199
transform 1 0 2400 0 -1 170
box -8 -3 16 105
use FILL  FILL_5170
timestamp 1711653199
transform 1 0 2360 0 -1 170
box -8 -3 16 105
use FILL  FILL_5171
timestamp 1711653199
transform 1 0 2352 0 -1 170
box -8 -3 16 105
use FILL  FILL_5172
timestamp 1711653199
transform 1 0 2312 0 -1 170
box -8 -3 16 105
use FILL  FILL_5173
timestamp 1711653199
transform 1 0 2304 0 -1 170
box -8 -3 16 105
use FILL  FILL_5174
timestamp 1711653199
transform 1 0 2296 0 -1 170
box -8 -3 16 105
use FILL  FILL_5175
timestamp 1711653199
transform 1 0 2288 0 -1 170
box -8 -3 16 105
use FILL  FILL_5176
timestamp 1711653199
transform 1 0 2280 0 -1 170
box -8 -3 16 105
use FILL  FILL_5177
timestamp 1711653199
transform 1 0 2272 0 -1 170
box -8 -3 16 105
use FILL  FILL_5178
timestamp 1711653199
transform 1 0 2216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5179
timestamp 1711653199
transform 1 0 2208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5180
timestamp 1711653199
transform 1 0 2200 0 -1 170
box -8 -3 16 105
use FILL  FILL_5181
timestamp 1711653199
transform 1 0 2192 0 -1 170
box -8 -3 16 105
use FILL  FILL_5182
timestamp 1711653199
transform 1 0 2184 0 -1 170
box -8 -3 16 105
use FILL  FILL_5183
timestamp 1711653199
transform 1 0 2176 0 -1 170
box -8 -3 16 105
use FILL  FILL_5184
timestamp 1711653199
transform 1 0 2152 0 -1 170
box -8 -3 16 105
use FILL  FILL_5185
timestamp 1711653199
transform 1 0 2104 0 -1 170
box -8 -3 16 105
use FILL  FILL_5186
timestamp 1711653199
transform 1 0 2096 0 -1 170
box -8 -3 16 105
use FILL  FILL_5187
timestamp 1711653199
transform 1 0 2088 0 -1 170
box -8 -3 16 105
use FILL  FILL_5188
timestamp 1711653199
transform 1 0 2080 0 -1 170
box -8 -3 16 105
use FILL  FILL_5189
timestamp 1711653199
transform 1 0 2072 0 -1 170
box -8 -3 16 105
use FILL  FILL_5190
timestamp 1711653199
transform 1 0 2064 0 -1 170
box -8 -3 16 105
use FILL  FILL_5191
timestamp 1711653199
transform 1 0 2016 0 -1 170
box -8 -3 16 105
use FILL  FILL_5192
timestamp 1711653199
transform 1 0 2008 0 -1 170
box -8 -3 16 105
use FILL  FILL_5193
timestamp 1711653199
transform 1 0 2000 0 -1 170
box -8 -3 16 105
use FILL  FILL_5194
timestamp 1711653199
transform 1 0 1992 0 -1 170
box -8 -3 16 105
use FILL  FILL_5195
timestamp 1711653199
transform 1 0 1984 0 -1 170
box -8 -3 16 105
use FILL  FILL_5196
timestamp 1711653199
transform 1 0 1944 0 -1 170
box -8 -3 16 105
use FILL  FILL_5197
timestamp 1711653199
transform 1 0 1936 0 -1 170
box -8 -3 16 105
use FILL  FILL_5198
timestamp 1711653199
transform 1 0 1928 0 -1 170
box -8 -3 16 105
use FILL  FILL_5199
timestamp 1711653199
transform 1 0 1888 0 -1 170
box -8 -3 16 105
use FILL  FILL_5200
timestamp 1711653199
transform 1 0 1880 0 -1 170
box -8 -3 16 105
use FILL  FILL_5201
timestamp 1711653199
transform 1 0 1872 0 -1 170
box -8 -3 16 105
use FILL  FILL_5202
timestamp 1711653199
transform 1 0 1864 0 -1 170
box -8 -3 16 105
use FILL  FILL_5203
timestamp 1711653199
transform 1 0 1856 0 -1 170
box -8 -3 16 105
use FILL  FILL_5204
timestamp 1711653199
transform 1 0 1848 0 -1 170
box -8 -3 16 105
use FILL  FILL_5205
timestamp 1711653199
transform 1 0 1840 0 -1 170
box -8 -3 16 105
use FILL  FILL_5206
timestamp 1711653199
transform 1 0 1792 0 -1 170
box -8 -3 16 105
use FILL  FILL_5207
timestamp 1711653199
transform 1 0 1784 0 -1 170
box -8 -3 16 105
use FILL  FILL_5208
timestamp 1711653199
transform 1 0 1776 0 -1 170
box -8 -3 16 105
use FILL  FILL_5209
timestamp 1711653199
transform 1 0 1768 0 -1 170
box -8 -3 16 105
use FILL  FILL_5210
timestamp 1711653199
transform 1 0 1760 0 -1 170
box -8 -3 16 105
use FILL  FILL_5211
timestamp 1711653199
transform 1 0 1752 0 -1 170
box -8 -3 16 105
use FILL  FILL_5212
timestamp 1711653199
transform 1 0 1720 0 -1 170
box -8 -3 16 105
use FILL  FILL_5213
timestamp 1711653199
transform 1 0 1712 0 -1 170
box -8 -3 16 105
use FILL  FILL_5214
timestamp 1711653199
transform 1 0 1680 0 -1 170
box -8 -3 16 105
use FILL  FILL_5215
timestamp 1711653199
transform 1 0 1672 0 -1 170
box -8 -3 16 105
use FILL  FILL_5216
timestamp 1711653199
transform 1 0 1664 0 -1 170
box -8 -3 16 105
use FILL  FILL_5217
timestamp 1711653199
transform 1 0 1656 0 -1 170
box -8 -3 16 105
use FILL  FILL_5218
timestamp 1711653199
transform 1 0 1648 0 -1 170
box -8 -3 16 105
use FILL  FILL_5219
timestamp 1711653199
transform 1 0 1640 0 -1 170
box -8 -3 16 105
use FILL  FILL_5220
timestamp 1711653199
transform 1 0 1600 0 -1 170
box -8 -3 16 105
use FILL  FILL_5221
timestamp 1711653199
transform 1 0 1592 0 -1 170
box -8 -3 16 105
use FILL  FILL_5222
timestamp 1711653199
transform 1 0 1584 0 -1 170
box -8 -3 16 105
use FILL  FILL_5223
timestamp 1711653199
transform 1 0 1576 0 -1 170
box -8 -3 16 105
use FILL  FILL_5224
timestamp 1711653199
transform 1 0 1568 0 -1 170
box -8 -3 16 105
use FILL  FILL_5225
timestamp 1711653199
transform 1 0 1528 0 -1 170
box -8 -3 16 105
use FILL  FILL_5226
timestamp 1711653199
transform 1 0 1520 0 -1 170
box -8 -3 16 105
use FILL  FILL_5227
timestamp 1711653199
transform 1 0 1512 0 -1 170
box -8 -3 16 105
use FILL  FILL_5228
timestamp 1711653199
transform 1 0 1504 0 -1 170
box -8 -3 16 105
use FILL  FILL_5229
timestamp 1711653199
transform 1 0 1496 0 -1 170
box -8 -3 16 105
use FILL  FILL_5230
timestamp 1711653199
transform 1 0 1488 0 -1 170
box -8 -3 16 105
use FILL  FILL_5231
timestamp 1711653199
transform 1 0 1448 0 -1 170
box -8 -3 16 105
use FILL  FILL_5232
timestamp 1711653199
transform 1 0 1440 0 -1 170
box -8 -3 16 105
use FILL  FILL_5233
timestamp 1711653199
transform 1 0 1432 0 -1 170
box -8 -3 16 105
use FILL  FILL_5234
timestamp 1711653199
transform 1 0 1424 0 -1 170
box -8 -3 16 105
use FILL  FILL_5235
timestamp 1711653199
transform 1 0 1416 0 -1 170
box -8 -3 16 105
use FILL  FILL_5236
timestamp 1711653199
transform 1 0 1384 0 -1 170
box -8 -3 16 105
use FILL  FILL_5237
timestamp 1711653199
transform 1 0 1376 0 -1 170
box -8 -3 16 105
use FILL  FILL_5238
timestamp 1711653199
transform 1 0 1368 0 -1 170
box -8 -3 16 105
use FILL  FILL_5239
timestamp 1711653199
transform 1 0 1360 0 -1 170
box -8 -3 16 105
use FILL  FILL_5240
timestamp 1711653199
transform 1 0 1312 0 -1 170
box -8 -3 16 105
use FILL  FILL_5241
timestamp 1711653199
transform 1 0 1304 0 -1 170
box -8 -3 16 105
use FILL  FILL_5242
timestamp 1711653199
transform 1 0 1296 0 -1 170
box -8 -3 16 105
use FILL  FILL_5243
timestamp 1711653199
transform 1 0 1288 0 -1 170
box -8 -3 16 105
use FILL  FILL_5244
timestamp 1711653199
transform 1 0 1280 0 -1 170
box -8 -3 16 105
use FILL  FILL_5245
timestamp 1711653199
transform 1 0 1272 0 -1 170
box -8 -3 16 105
use FILL  FILL_5246
timestamp 1711653199
transform 1 0 1224 0 -1 170
box -8 -3 16 105
use FILL  FILL_5247
timestamp 1711653199
transform 1 0 1216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5248
timestamp 1711653199
transform 1 0 1208 0 -1 170
box -8 -3 16 105
use FILL  FILL_5249
timestamp 1711653199
transform 1 0 1200 0 -1 170
box -8 -3 16 105
use FILL  FILL_5250
timestamp 1711653199
transform 1 0 1192 0 -1 170
box -8 -3 16 105
use FILL  FILL_5251
timestamp 1711653199
transform 1 0 1144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5252
timestamp 1711653199
transform 1 0 1136 0 -1 170
box -8 -3 16 105
use FILL  FILL_5253
timestamp 1711653199
transform 1 0 1128 0 -1 170
box -8 -3 16 105
use FILL  FILL_5254
timestamp 1711653199
transform 1 0 1120 0 -1 170
box -8 -3 16 105
use FILL  FILL_5255
timestamp 1711653199
transform 1 0 1112 0 -1 170
box -8 -3 16 105
use FILL  FILL_5256
timestamp 1711653199
transform 1 0 1104 0 -1 170
box -8 -3 16 105
use FILL  FILL_5257
timestamp 1711653199
transform 1 0 1064 0 -1 170
box -8 -3 16 105
use FILL  FILL_5258
timestamp 1711653199
transform 1 0 1056 0 -1 170
box -8 -3 16 105
use FILL  FILL_5259
timestamp 1711653199
transform 1 0 1016 0 -1 170
box -8 -3 16 105
use FILL  FILL_5260
timestamp 1711653199
transform 1 0 1008 0 -1 170
box -8 -3 16 105
use FILL  FILL_5261
timestamp 1711653199
transform 1 0 1000 0 -1 170
box -8 -3 16 105
use FILL  FILL_5262
timestamp 1711653199
transform 1 0 992 0 -1 170
box -8 -3 16 105
use FILL  FILL_5263
timestamp 1711653199
transform 1 0 984 0 -1 170
box -8 -3 16 105
use FILL  FILL_5264
timestamp 1711653199
transform 1 0 976 0 -1 170
box -8 -3 16 105
use FILL  FILL_5265
timestamp 1711653199
transform 1 0 944 0 -1 170
box -8 -3 16 105
use FILL  FILL_5266
timestamp 1711653199
transform 1 0 912 0 -1 170
box -8 -3 16 105
use FILL  FILL_5267
timestamp 1711653199
transform 1 0 904 0 -1 170
box -8 -3 16 105
use FILL  FILL_5268
timestamp 1711653199
transform 1 0 896 0 -1 170
box -8 -3 16 105
use FILL  FILL_5269
timestamp 1711653199
transform 1 0 888 0 -1 170
box -8 -3 16 105
use FILL  FILL_5270
timestamp 1711653199
transform 1 0 880 0 -1 170
box -8 -3 16 105
use FILL  FILL_5271
timestamp 1711653199
transform 1 0 872 0 -1 170
box -8 -3 16 105
use FILL  FILL_5272
timestamp 1711653199
transform 1 0 824 0 -1 170
box -8 -3 16 105
use FILL  FILL_5273
timestamp 1711653199
transform 1 0 816 0 -1 170
box -8 -3 16 105
use FILL  FILL_5274
timestamp 1711653199
transform 1 0 808 0 -1 170
box -8 -3 16 105
use FILL  FILL_5275
timestamp 1711653199
transform 1 0 800 0 -1 170
box -8 -3 16 105
use FILL  FILL_5276
timestamp 1711653199
transform 1 0 792 0 -1 170
box -8 -3 16 105
use FILL  FILL_5277
timestamp 1711653199
transform 1 0 784 0 -1 170
box -8 -3 16 105
use FILL  FILL_5278
timestamp 1711653199
transform 1 0 736 0 -1 170
box -8 -3 16 105
use FILL  FILL_5279
timestamp 1711653199
transform 1 0 728 0 -1 170
box -8 -3 16 105
use FILL  FILL_5280
timestamp 1711653199
transform 1 0 720 0 -1 170
box -8 -3 16 105
use FILL  FILL_5281
timestamp 1711653199
transform 1 0 712 0 -1 170
box -8 -3 16 105
use FILL  FILL_5282
timestamp 1711653199
transform 1 0 704 0 -1 170
box -8 -3 16 105
use FILL  FILL_5283
timestamp 1711653199
transform 1 0 672 0 -1 170
box -8 -3 16 105
use FILL  FILL_5284
timestamp 1711653199
transform 1 0 664 0 -1 170
box -8 -3 16 105
use FILL  FILL_5285
timestamp 1711653199
transform 1 0 656 0 -1 170
box -8 -3 16 105
use FILL  FILL_5286
timestamp 1711653199
transform 1 0 648 0 -1 170
box -8 -3 16 105
use FILL  FILL_5287
timestamp 1711653199
transform 1 0 640 0 -1 170
box -8 -3 16 105
use FILL  FILL_5288
timestamp 1711653199
transform 1 0 592 0 -1 170
box -8 -3 16 105
use FILL  FILL_5289
timestamp 1711653199
transform 1 0 584 0 -1 170
box -8 -3 16 105
use FILL  FILL_5290
timestamp 1711653199
transform 1 0 576 0 -1 170
box -8 -3 16 105
use FILL  FILL_5291
timestamp 1711653199
transform 1 0 568 0 -1 170
box -8 -3 16 105
use FILL  FILL_5292
timestamp 1711653199
transform 1 0 560 0 -1 170
box -8 -3 16 105
use FILL  FILL_5293
timestamp 1711653199
transform 1 0 528 0 -1 170
box -8 -3 16 105
use FILL  FILL_5294
timestamp 1711653199
transform 1 0 520 0 -1 170
box -8 -3 16 105
use FILL  FILL_5295
timestamp 1711653199
transform 1 0 512 0 -1 170
box -8 -3 16 105
use FILL  FILL_5296
timestamp 1711653199
transform 1 0 488 0 -1 170
box -8 -3 16 105
use FILL  FILL_5297
timestamp 1711653199
transform 1 0 480 0 -1 170
box -8 -3 16 105
use FILL  FILL_5298
timestamp 1711653199
transform 1 0 472 0 -1 170
box -8 -3 16 105
use FILL  FILL_5299
timestamp 1711653199
transform 1 0 424 0 -1 170
box -8 -3 16 105
use FILL  FILL_5300
timestamp 1711653199
transform 1 0 416 0 -1 170
box -8 -3 16 105
use FILL  FILL_5301
timestamp 1711653199
transform 1 0 408 0 -1 170
box -8 -3 16 105
use FILL  FILL_5302
timestamp 1711653199
transform 1 0 400 0 -1 170
box -8 -3 16 105
use FILL  FILL_5303
timestamp 1711653199
transform 1 0 392 0 -1 170
box -8 -3 16 105
use FILL  FILL_5304
timestamp 1711653199
transform 1 0 384 0 -1 170
box -8 -3 16 105
use FILL  FILL_5305
timestamp 1711653199
transform 1 0 336 0 -1 170
box -8 -3 16 105
use FILL  FILL_5306
timestamp 1711653199
transform 1 0 328 0 -1 170
box -8 -3 16 105
use FILL  FILL_5307
timestamp 1711653199
transform 1 0 320 0 -1 170
box -8 -3 16 105
use FILL  FILL_5308
timestamp 1711653199
transform 1 0 312 0 -1 170
box -8 -3 16 105
use FILL  FILL_5309
timestamp 1711653199
transform 1 0 304 0 -1 170
box -8 -3 16 105
use FILL  FILL_5310
timestamp 1711653199
transform 1 0 256 0 -1 170
box -8 -3 16 105
use FILL  FILL_5311
timestamp 1711653199
transform 1 0 248 0 -1 170
box -8 -3 16 105
use FILL  FILL_5312
timestamp 1711653199
transform 1 0 240 0 -1 170
box -8 -3 16 105
use FILL  FILL_5313
timestamp 1711653199
transform 1 0 232 0 -1 170
box -8 -3 16 105
use FILL  FILL_5314
timestamp 1711653199
transform 1 0 224 0 -1 170
box -8 -3 16 105
use FILL  FILL_5315
timestamp 1711653199
transform 1 0 216 0 -1 170
box -8 -3 16 105
use FILL  FILL_5316
timestamp 1711653199
transform 1 0 168 0 -1 170
box -8 -3 16 105
use FILL  FILL_5317
timestamp 1711653199
transform 1 0 160 0 -1 170
box -8 -3 16 105
use FILL  FILL_5318
timestamp 1711653199
transform 1 0 152 0 -1 170
box -8 -3 16 105
use FILL  FILL_5319
timestamp 1711653199
transform 1 0 144 0 -1 170
box -8 -3 16 105
use FILL  FILL_5320
timestamp 1711653199
transform 1 0 136 0 -1 170
box -8 -3 16 105
use FILL  FILL_5321
timestamp 1711653199
transform 1 0 104 0 -1 170
box -8 -3 16 105
use FILL  FILL_5322
timestamp 1711653199
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_5323
timestamp 1711653199
transform 1 0 88 0 -1 170
box -8 -3 16 105
use FILL  FILL_5324
timestamp 1711653199
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_5325
timestamp 1711653199
transform 1 0 72 0 -1 170
box -8 -3 16 105
use HAX1  HAX1_0
timestamp 1711653199
transform 1 0 2712 0 -1 2770
box -5 -3 84 105
use HAX1  HAX1_1
timestamp 1711653199
transform 1 0 2808 0 -1 2770
box -5 -3 84 105
use HAX1  HAX1_2
timestamp 1711653199
transform 1 0 2936 0 -1 2770
box -5 -3 84 105
use INVX2  INVX2_0
timestamp 1711653199
transform 1 0 3192 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_1
timestamp 1711653199
transform 1 0 2944 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_2
timestamp 1711653199
transform 1 0 3136 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_3
timestamp 1711653199
transform 1 0 1512 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_4
timestamp 1711653199
transform 1 0 2888 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_5
timestamp 1711653199
transform 1 0 2632 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_6
timestamp 1711653199
transform 1 0 1704 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_7
timestamp 1711653199
transform 1 0 2952 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_8
timestamp 1711653199
transform 1 0 2336 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_9
timestamp 1711653199
transform 1 0 2976 0 1 770
box -9 -3 26 105
use INVX2  INVX2_10
timestamp 1711653199
transform 1 0 2936 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_11
timestamp 1711653199
transform 1 0 512 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_12
timestamp 1711653199
transform 1 0 528 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_13
timestamp 1711653199
transform 1 0 2032 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_14
timestamp 1711653199
transform 1 0 664 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_15
timestamp 1711653199
transform 1 0 832 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_16
timestamp 1711653199
transform 1 0 2952 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_17
timestamp 1711653199
transform 1 0 2640 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_18
timestamp 1711653199
transform 1 0 2200 0 1 770
box -9 -3 26 105
use INVX2  INVX2_19
timestamp 1711653199
transform 1 0 248 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_20
timestamp 1711653199
transform 1 0 2944 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_21
timestamp 1711653199
transform 1 0 2696 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_22
timestamp 1711653199
transform 1 0 2632 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_23
timestamp 1711653199
transform 1 0 2128 0 1 970
box -9 -3 26 105
use INVX2  INVX2_24
timestamp 1711653199
transform 1 0 1656 0 1 570
box -9 -3 26 105
use INVX2  INVX2_25
timestamp 1711653199
transform 1 0 2256 0 1 570
box -9 -3 26 105
use INVX2  INVX2_26
timestamp 1711653199
transform 1 0 2600 0 1 770
box -9 -3 26 105
use INVX2  INVX2_27
timestamp 1711653199
transform 1 0 1000 0 1 370
box -9 -3 26 105
use INVX2  INVX2_28
timestamp 1711653199
transform 1 0 1312 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_29
timestamp 1711653199
transform 1 0 2152 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_30
timestamp 1711653199
transform 1 0 232 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_31
timestamp 1711653199
transform 1 0 1144 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_32
timestamp 1711653199
transform 1 0 2760 0 1 770
box -9 -3 26 105
use INVX2  INVX2_33
timestamp 1711653199
transform 1 0 2696 0 1 970
box -9 -3 26 105
use INVX2  INVX2_34
timestamp 1711653199
transform 1 0 2216 0 1 770
box -9 -3 26 105
use INVX2  INVX2_35
timestamp 1711653199
transform 1 0 2592 0 1 170
box -9 -3 26 105
use INVX2  INVX2_36
timestamp 1711653199
transform 1 0 2496 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_37
timestamp 1711653199
transform 1 0 2856 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_38
timestamp 1711653199
transform 1 0 2440 0 1 770
box -9 -3 26 105
use INVX2  INVX2_39
timestamp 1711653199
transform 1 0 1736 0 1 170
box -9 -3 26 105
use INVX2  INVX2_40
timestamp 1711653199
transform 1 0 1856 0 1 370
box -9 -3 26 105
use INVX2  INVX2_41
timestamp 1711653199
transform 1 0 2128 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_42
timestamp 1711653199
transform 1 0 2104 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_43
timestamp 1711653199
transform 1 0 2240 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_44
timestamp 1711653199
transform 1 0 2368 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_45
timestamp 1711653199
transform 1 0 1048 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_46
timestamp 1711653199
transform 1 0 736 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_47
timestamp 1711653199
transform 1 0 2304 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_48
timestamp 1711653199
transform 1 0 696 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_49
timestamp 1711653199
transform 1 0 2728 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_50
timestamp 1711653199
transform 1 0 1120 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_51
timestamp 1711653199
transform 1 0 296 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_52
timestamp 1711653199
transform 1 0 480 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_53
timestamp 1711653199
transform 1 0 2496 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_54
timestamp 1711653199
transform 1 0 2384 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_55
timestamp 1711653199
transform 1 0 1696 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_56
timestamp 1711653199
transform 1 0 1064 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_57
timestamp 1711653199
transform 1 0 1328 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_58
timestamp 1711653199
transform 1 0 2064 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_59
timestamp 1711653199
transform 1 0 2520 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_60
timestamp 1711653199
transform 1 0 1768 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_61
timestamp 1711653199
transform 1 0 2304 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_62
timestamp 1711653199
transform 1 0 672 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_63
timestamp 1711653199
transform 1 0 656 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_64
timestamp 1711653199
transform 1 0 2992 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_65
timestamp 1711653199
transform 1 0 1680 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_66
timestamp 1711653199
transform 1 0 1752 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_67
timestamp 1711653199
transform 1 0 568 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_68
timestamp 1711653199
transform 1 0 824 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_69
timestamp 1711653199
transform 1 0 2240 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_70
timestamp 1711653199
transform 1 0 2952 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_71
timestamp 1711653199
transform 1 0 1864 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_72
timestamp 1711653199
transform 1 0 1960 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_73
timestamp 1711653199
transform 1 0 400 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_74
timestamp 1711653199
transform 1 0 1496 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_75
timestamp 1711653199
transform 1 0 2920 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_76
timestamp 1711653199
transform 1 0 1904 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_77
timestamp 1711653199
transform 1 0 792 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_78
timestamp 1711653199
transform 1 0 624 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_79
timestamp 1711653199
transform 1 0 2864 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_80
timestamp 1711653199
transform 1 0 2168 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_81
timestamp 1711653199
transform 1 0 1208 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_82
timestamp 1711653199
transform 1 0 1992 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_83
timestamp 1711653199
transform 1 0 1808 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_84
timestamp 1711653199
transform 1 0 1608 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_85
timestamp 1711653199
transform 1 0 1368 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_86
timestamp 1711653199
transform 1 0 888 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_87
timestamp 1711653199
transform 1 0 672 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_88
timestamp 1711653199
transform 1 0 328 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_89
timestamp 1711653199
transform 1 0 512 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_90
timestamp 1711653199
transform 1 0 192 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_91
timestamp 1711653199
transform 1 0 200 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_92
timestamp 1711653199
transform 1 0 248 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_93
timestamp 1711653199
transform 1 0 184 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_94
timestamp 1711653199
transform 1 0 272 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_95
timestamp 1711653199
transform 1 0 312 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_96
timestamp 1711653199
transform 1 0 432 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_97
timestamp 1711653199
transform 1 0 728 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_98
timestamp 1711653199
transform 1 0 1120 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_99
timestamp 1711653199
transform 1 0 816 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_100
timestamp 1711653199
transform 1 0 984 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_101
timestamp 1711653199
transform 1 0 1264 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_102
timestamp 1711653199
transform 1 0 1480 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_103
timestamp 1711653199
transform 1 0 1680 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_104
timestamp 1711653199
transform 1 0 1616 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_105
timestamp 1711653199
transform 1 0 1848 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_106
timestamp 1711653199
transform 1 0 1912 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_107
timestamp 1711653199
transform 1 0 2256 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_108
timestamp 1711653199
transform 1 0 2176 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_109
timestamp 1711653199
transform 1 0 2464 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_110
timestamp 1711653199
transform 1 0 2424 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_111
timestamp 1711653199
transform 1 0 2016 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_112
timestamp 1711653199
transform 1 0 3160 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_113
timestamp 1711653199
transform 1 0 2704 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_114
timestamp 1711653199
transform 1 0 3296 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_115
timestamp 1711653199
transform 1 0 3064 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_116
timestamp 1711653199
transform 1 0 3136 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_117
timestamp 1711653199
transform 1 0 3120 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_118
timestamp 1711653199
transform 1 0 3360 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_119
timestamp 1711653199
transform 1 0 3360 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_120
timestamp 1711653199
transform 1 0 2736 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_121
timestamp 1711653199
transform 1 0 2768 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_122
timestamp 1711653199
transform 1 0 2864 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_123
timestamp 1711653199
transform 1 0 3184 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_124
timestamp 1711653199
transform 1 0 3224 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_125
timestamp 1711653199
transform 1 0 3232 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_126
timestamp 1711653199
transform 1 0 3056 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_127
timestamp 1711653199
transform 1 0 3016 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_128
timestamp 1711653199
transform 1 0 3216 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_129
timestamp 1711653199
transform 1 0 1128 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_130
timestamp 1711653199
transform 1 0 952 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_131
timestamp 1711653199
transform 1 0 936 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_132
timestamp 1711653199
transform 1 0 1096 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_133
timestamp 1711653199
transform 1 0 2160 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_134
timestamp 1711653199
transform 1 0 2440 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_135
timestamp 1711653199
transform 1 0 2480 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_136
timestamp 1711653199
transform 1 0 1232 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_137
timestamp 1711653199
transform 1 0 2984 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_138
timestamp 1711653199
transform 1 0 2912 0 1 170
box -9 -3 26 105
use INVX2  INVX2_139
timestamp 1711653199
transform 1 0 3088 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_140
timestamp 1711653199
transform 1 0 3024 0 1 370
box -9 -3 26 105
use INVX2  INVX2_141
timestamp 1711653199
transform 1 0 3056 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_142
timestamp 1711653199
transform 1 0 2976 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_143
timestamp 1711653199
transform 1 0 1896 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_144
timestamp 1711653199
transform 1 0 3320 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_145
timestamp 1711653199
transform 1 0 3304 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_146
timestamp 1711653199
transform 1 0 2152 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_147
timestamp 1711653199
transform 1 0 3360 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_148
timestamp 1711653199
transform 1 0 3336 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_149
timestamp 1711653199
transform 1 0 3368 0 1 570
box -9 -3 26 105
use INVX2  INVX2_150
timestamp 1711653199
transform 1 0 2672 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_151
timestamp 1711653199
transform 1 0 1440 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_152
timestamp 1711653199
transform 1 0 2752 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_153
timestamp 1711653199
transform 1 0 2632 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_154
timestamp 1711653199
transform 1 0 2656 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_155
timestamp 1711653199
transform 1 0 2848 0 1 170
box -9 -3 26 105
use INVX2  INVX2_156
timestamp 1711653199
transform 1 0 2736 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_157
timestamp 1711653199
transform 1 0 2744 0 1 770
box -9 -3 26 105
use INVX2  INVX2_158
timestamp 1711653199
transform 1 0 2128 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_159
timestamp 1711653199
transform 1 0 2048 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_160
timestamp 1711653199
transform 1 0 2080 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_161
timestamp 1711653199
transform 1 0 2136 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_162
timestamp 1711653199
transform 1 0 1752 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_163
timestamp 1711653199
transform 1 0 1648 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_164
timestamp 1711653199
transform 1 0 2040 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_165
timestamp 1711653199
transform 1 0 2520 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_166
timestamp 1711653199
transform 1 0 2392 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_167
timestamp 1711653199
transform 1 0 1704 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_168
timestamp 1711653199
transform 1 0 2560 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_169
timestamp 1711653199
transform 1 0 2192 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_170
timestamp 1711653199
transform 1 0 2600 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_171
timestamp 1711653199
transform 1 0 2328 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_172
timestamp 1711653199
transform 1 0 1968 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_173
timestamp 1711653199
transform 1 0 1232 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_174
timestamp 1711653199
transform 1 0 1952 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_175
timestamp 1711653199
transform 1 0 2352 0 1 770
box -9 -3 26 105
use INVX2  INVX2_176
timestamp 1711653199
transform 1 0 2360 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_177
timestamp 1711653199
transform 1 0 2560 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_178
timestamp 1711653199
transform 1 0 2120 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_179
timestamp 1711653199
transform 1 0 1728 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_180
timestamp 1711653199
transform 1 0 2080 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_181
timestamp 1711653199
transform 1 0 2040 0 1 770
box -9 -3 26 105
use INVX2  INVX2_182
timestamp 1711653199
transform 1 0 2056 0 1 970
box -9 -3 26 105
use INVX2  INVX2_183
timestamp 1711653199
transform 1 0 1728 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_184
timestamp 1711653199
transform 1 0 1800 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_185
timestamp 1711653199
transform 1 0 1304 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_186
timestamp 1711653199
transform 1 0 1960 0 1 970
box -9 -3 26 105
use INVX2  INVX2_187
timestamp 1711653199
transform 1 0 1936 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_188
timestamp 1711653199
transform 1 0 1528 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_189
timestamp 1711653199
transform 1 0 1176 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_190
timestamp 1711653199
transform 1 0 1832 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_191
timestamp 1711653199
transform 1 0 2480 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_192
timestamp 1711653199
transform 1 0 1832 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_193
timestamp 1711653199
transform 1 0 1496 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_194
timestamp 1711653199
transform 1 0 992 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_195
timestamp 1711653199
transform 1 0 1136 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_196
timestamp 1711653199
transform 1 0 1936 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_197
timestamp 1711653199
transform 1 0 2200 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_198
timestamp 1711653199
transform 1 0 1008 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_199
timestamp 1711653199
transform 1 0 704 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_200
timestamp 1711653199
transform 1 0 672 0 1 170
box -9 -3 26 105
use INVX2  INVX2_201
timestamp 1711653199
transform 1 0 624 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_202
timestamp 1711653199
transform 1 0 1128 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_203
timestamp 1711653199
transform 1 0 248 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_204
timestamp 1711653199
transform 1 0 328 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_205
timestamp 1711653199
transform 1 0 1144 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_206
timestamp 1711653199
transform 1 0 264 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_207
timestamp 1711653199
transform 1 0 168 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_208
timestamp 1711653199
transform 1 0 88 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_209
timestamp 1711653199
transform 1 0 88 0 1 970
box -9 -3 26 105
use INVX2  INVX2_210
timestamp 1711653199
transform 1 0 88 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_211
timestamp 1711653199
transform 1 0 1120 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_212
timestamp 1711653199
transform 1 0 896 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_213
timestamp 1711653199
transform 1 0 984 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_214
timestamp 1711653199
transform 1 0 1232 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_215
timestamp 1711653199
transform 1 0 408 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_216
timestamp 1711653199
transform 1 0 80 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_217
timestamp 1711653199
transform 1 0 2136 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_218
timestamp 1711653199
transform 1 0 880 0 1 970
box -9 -3 26 105
use INVX2  INVX2_219
timestamp 1711653199
transform 1 0 512 0 1 970
box -9 -3 26 105
use INVX2  INVX2_220
timestamp 1711653199
transform 1 0 512 0 1 370
box -9 -3 26 105
use INVX2  INVX2_221
timestamp 1711653199
transform 1 0 872 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_222
timestamp 1711653199
transform 1 0 520 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_223
timestamp 1711653199
transform 1 0 720 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_224
timestamp 1711653199
transform 1 0 752 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_225
timestamp 1711653199
transform 1 0 680 0 1 970
box -9 -3 26 105
use INVX2  INVX2_226
timestamp 1711653199
transform 1 0 688 0 1 770
box -9 -3 26 105
use INVX2  INVX2_227
timestamp 1711653199
transform 1 0 400 0 1 770
box -9 -3 26 105
use INVX2  INVX2_228
timestamp 1711653199
transform 1 0 736 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_229
timestamp 1711653199
transform 1 0 848 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_230
timestamp 1711653199
transform 1 0 976 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_231
timestamp 1711653199
transform 1 0 616 0 1 570
box -9 -3 26 105
use INVX2  INVX2_232
timestamp 1711653199
transform 1 0 752 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_233
timestamp 1711653199
transform 1 0 1104 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_234
timestamp 1711653199
transform 1 0 2344 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_235
timestamp 1711653199
transform 1 0 1752 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_236
timestamp 1711653199
transform 1 0 984 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_237
timestamp 1711653199
transform 1 0 880 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_238
timestamp 1711653199
transform 1 0 928 0 -1 1570
box -9 -3 26 105
use INVX2  INVX2_239
timestamp 1711653199
transform 1 0 880 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_240
timestamp 1711653199
transform 1 0 776 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_241
timestamp 1711653199
transform 1 0 760 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_242
timestamp 1711653199
transform 1 0 432 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_243
timestamp 1711653199
transform 1 0 496 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_244
timestamp 1711653199
transform 1 0 440 0 1 370
box -9 -3 26 105
use INVX2  INVX2_245
timestamp 1711653199
transform 1 0 680 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_246
timestamp 1711653199
transform 1 0 88 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_247
timestamp 1711653199
transform 1 0 232 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_248
timestamp 1711653199
transform 1 0 816 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_249
timestamp 1711653199
transform 1 0 896 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_250
timestamp 1711653199
transform 1 0 1040 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_251
timestamp 1711653199
transform 1 0 1552 0 1 170
box -9 -3 26 105
use INVX2  INVX2_252
timestamp 1711653199
transform 1 0 880 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_253
timestamp 1711653199
transform 1 0 936 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_254
timestamp 1711653199
transform 1 0 1032 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_255
timestamp 1711653199
transform 1 0 1088 0 1 170
box -9 -3 26 105
use INVX2  INVX2_256
timestamp 1711653199
transform 1 0 1320 0 1 370
box -9 -3 26 105
use INVX2  INVX2_257
timestamp 1711653199
transform 1 0 1144 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_258
timestamp 1711653199
transform 1 0 936 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_259
timestamp 1711653199
transform 1 0 1504 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_260
timestamp 1711653199
transform 1 0 1104 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_261
timestamp 1711653199
transform 1 0 1520 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_262
timestamp 1711653199
transform 1 0 2216 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_263
timestamp 1711653199
transform 1 0 1232 0 1 970
box -9 -3 26 105
use INVX2  INVX2_264
timestamp 1711653199
transform 1 0 1256 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_265
timestamp 1711653199
transform 1 0 1184 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_266
timestamp 1711653199
transform 1 0 920 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_267
timestamp 1711653199
transform 1 0 2264 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_268
timestamp 1711653199
transform 1 0 1976 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_269
timestamp 1711653199
transform 1 0 2960 0 -1 1970
box -9 -3 26 105
use INVX2  INVX2_270
timestamp 1711653199
transform 1 0 3064 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_271
timestamp 1711653199
transform 1 0 2064 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_272
timestamp 1711653199
transform 1 0 3344 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_273
timestamp 1711653199
transform 1 0 3288 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_274
timestamp 1711653199
transform 1 0 3272 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_275
timestamp 1711653199
transform 1 0 3368 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_276
timestamp 1711653199
transform 1 0 3344 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_277
timestamp 1711653199
transform 1 0 3336 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_278
timestamp 1711653199
transform 1 0 3360 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_279
timestamp 1711653199
transform 1 0 3008 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_280
timestamp 1711653199
transform 1 0 2952 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_281
timestamp 1711653199
transform 1 0 2400 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_282
timestamp 1711653199
transform 1 0 2608 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_283
timestamp 1711653199
transform 1 0 2464 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_284
timestamp 1711653199
transform 1 0 2704 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_285
timestamp 1711653199
transform 1 0 1904 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_286
timestamp 1711653199
transform 1 0 280 0 1 370
box -9 -3 26 105
use INVX2  INVX2_287
timestamp 1711653199
transform 1 0 2240 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_288
timestamp 1711653199
transform 1 0 1144 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_289
timestamp 1711653199
transform 1 0 2352 0 1 970
box -9 -3 26 105
use INVX2  INVX2_290
timestamp 1711653199
transform 1 0 2568 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_291
timestamp 1711653199
transform 1 0 944 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_292
timestamp 1711653199
transform 1 0 3224 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_293
timestamp 1711653199
transform 1 0 2480 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_294
timestamp 1711653199
transform 1 0 3040 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_295
timestamp 1711653199
transform 1 0 2600 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_296
timestamp 1711653199
transform 1 0 3152 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_297
timestamp 1711653199
transform 1 0 2840 0 1 570
box -9 -3 26 105
use INVX2  INVX2_298
timestamp 1711653199
transform 1 0 2976 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_299
timestamp 1711653199
transform 1 0 872 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_300
timestamp 1711653199
transform 1 0 320 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_301
timestamp 1711653199
transform 1 0 1520 0 1 2170
box -9 -3 26 105
use INVX2  INVX2_302
timestamp 1711653199
transform 1 0 2320 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_303
timestamp 1711653199
transform 1 0 2808 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_304
timestamp 1711653199
transform 1 0 2800 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_305
timestamp 1711653199
transform 1 0 2200 0 1 970
box -9 -3 26 105
use INVX2  INVX2_306
timestamp 1711653199
transform 1 0 3088 0 1 970
box -9 -3 26 105
use INVX2  INVX2_307
timestamp 1711653199
transform 1 0 3056 0 1 570
box -9 -3 26 105
use INVX2  INVX2_308
timestamp 1711653199
transform 1 0 2912 0 -1 1770
box -9 -3 26 105
use INVX2  INVX2_309
timestamp 1711653199
transform 1 0 3160 0 1 1570
box -9 -3 26 105
use INVX2  INVX2_310
timestamp 1711653199
transform 1 0 1104 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_311
timestamp 1711653199
transform 1 0 2864 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_312
timestamp 1711653199
transform 1 0 2808 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_313
timestamp 1711653199
transform 1 0 2720 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_314
timestamp 1711653199
transform 1 0 2736 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_315
timestamp 1711653199
transform 1 0 240 0 1 370
box -9 -3 26 105
use INVX2  INVX2_316
timestamp 1711653199
transform 1 0 2800 0 1 370
box -9 -3 26 105
use INVX2  INVX2_317
timestamp 1711653199
transform 1 0 1944 0 1 370
box -9 -3 26 105
use INVX2  INVX2_318
timestamp 1711653199
transform 1 0 2896 0 1 170
box -9 -3 26 105
use INVX2  INVX2_319
timestamp 1711653199
transform 1 0 2560 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_320
timestamp 1711653199
transform 1 0 2040 0 1 1970
box -9 -3 26 105
use INVX2  INVX2_321
timestamp 1711653199
transform 1 0 2912 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_322
timestamp 1711653199
transform 1 0 2360 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_323
timestamp 1711653199
transform 1 0 2152 0 -1 2770
box -9 -3 26 105
use INVX2  INVX2_324
timestamp 1711653199
transform 1 0 2304 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_325
timestamp 1711653199
transform 1 0 2720 0 -1 170
box -9 -3 26 105
use INVX2  INVX2_326
timestamp 1711653199
transform 1 0 2656 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_327
timestamp 1711653199
transform 1 0 2592 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_328
timestamp 1711653199
transform 1 0 2408 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_329
timestamp 1711653199
transform 1 0 3040 0 1 570
box -9 -3 26 105
use INVX2  INVX2_330
timestamp 1711653199
transform 1 0 1712 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_331
timestamp 1711653199
transform 1 0 1664 0 1 970
box -9 -3 26 105
use INVX2  INVX2_332
timestamp 1711653199
transform 1 0 1776 0 1 970
box -9 -3 26 105
use INVX2  INVX2_333
timestamp 1711653199
transform 1 0 3144 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_334
timestamp 1711653199
transform 1 0 3192 0 -1 2570
box -9 -3 26 105
use INVX2  INVX2_335
timestamp 1711653199
transform 1 0 3152 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_336
timestamp 1711653199
transform 1 0 3344 0 1 1770
box -9 -3 26 105
use INVX2  INVX2_337
timestamp 1711653199
transform 1 0 3008 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_338
timestamp 1711653199
transform 1 0 3120 0 1 2770
box -9 -3 26 105
use M2_M1  M2_M1_0
timestamp 1711653199
transform 1 0 2964 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1711653199
transform 1 0 2820 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1711653199
transform 1 0 2836 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1711653199
transform 1 0 2724 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1711653199
transform 1 0 2740 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_5
timestamp 1711653199
transform 1 0 2652 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1711653199
transform 1 0 2692 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1711653199
transform 1 0 2420 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1711653199
transform 1 0 2388 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_9
timestamp 1711653199
transform 1 0 2340 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1711653199
transform 1 0 2308 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_11
timestamp 1711653199
transform 1 0 2260 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1711653199
transform 1 0 2548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1711653199
transform 1 0 2396 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_14
timestamp 1711653199
transform 1 0 2324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1711653199
transform 1 0 2324 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1711653199
transform 1 0 2292 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1711653199
transform 1 0 2292 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1711653199
transform 1 0 2540 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1711653199
transform 1 0 2420 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1711653199
transform 1 0 2308 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_21
timestamp 1711653199
transform 1 0 2260 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1711653199
transform 1 0 2244 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1711653199
transform 1 0 2244 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1711653199
transform 1 0 2580 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_25
timestamp 1711653199
transform 1 0 2524 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1711653199
transform 1 0 2124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1711653199
transform 1 0 2108 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1711653199
transform 1 0 2644 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1711653199
transform 1 0 2548 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1711653199
transform 1 0 2124 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1711653199
transform 1 0 2076 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1711653199
transform 1 0 3348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1711653199
transform 1 0 3332 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1711653199
transform 1 0 3276 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1711653199
transform 1 0 2932 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1711653199
transform 1 0 2828 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1711653199
transform 1 0 2332 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1711653199
transform 1 0 2300 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1711653199
transform 1 0 1956 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1711653199
transform 1 0 948 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1711653199
transform 1 0 828 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1711653199
transform 1 0 828 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_43
timestamp 1711653199
transform 1 0 644 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1711653199
transform 1 0 604 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1711653199
transform 1 0 420 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1711653199
transform 1 0 324 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1711653199
transform 1 0 268 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1711653199
transform 1 0 220 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1711653199
transform 1 0 84 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1711653199
transform 1 0 3060 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_51
timestamp 1711653199
transform 1 0 2916 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_52
timestamp 1711653199
transform 1 0 2884 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1711653199
transform 1 0 2820 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1711653199
transform 1 0 3116 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1711653199
transform 1 0 3004 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1711653199
transform 1 0 2980 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1711653199
transform 1 0 2924 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1711653199
transform 1 0 2828 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1711653199
transform 1 0 2828 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1711653199
transform 1 0 3012 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1711653199
transform 1 0 2956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1711653199
transform 1 0 2956 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1711653199
transform 1 0 2892 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1711653199
transform 1 0 2892 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_65
timestamp 1711653199
transform 1 0 2836 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1711653199
transform 1 0 2772 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1711653199
transform 1 0 2740 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1711653199
transform 1 0 2708 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1711653199
transform 1 0 2884 0 1 1645
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1711653199
transform 1 0 2860 0 1 1645
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1711653199
transform 1 0 2804 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1711653199
transform 1 0 2740 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1711653199
transform 1 0 2716 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1711653199
transform 1 0 2692 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1711653199
transform 1 0 2660 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1711653199
transform 1 0 2636 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1711653199
transform 1 0 2724 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1711653199
transform 1 0 2692 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1711653199
transform 1 0 2692 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1711653199
transform 1 0 2652 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1711653199
transform 1 0 2596 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1711653199
transform 1 0 2572 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1711653199
transform 1 0 3372 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1711653199
transform 1 0 3204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1711653199
transform 1 0 3124 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1711653199
transform 1 0 3116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1711653199
transform 1 0 3068 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1711653199
transform 1 0 3300 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1711653199
transform 1 0 3196 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1711653199
transform 1 0 3108 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1711653199
transform 1 0 2076 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1711653199
transform 1 0 2020 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1711653199
transform 1 0 2572 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1711653199
transform 1 0 2468 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1711653199
transform 1 0 2300 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1711653199
transform 1 0 2260 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1711653199
transform 1 0 2620 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1711653199
transform 1 0 2604 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1711653199
transform 1 0 2508 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1711653199
transform 1 0 2524 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_101
timestamp 1711653199
transform 1 0 2476 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1711653199
transform 1 0 2380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1711653199
transform 1 0 1980 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1711653199
transform 1 0 1916 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1711653199
transform 1 0 1740 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1711653199
transform 1 0 1684 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1711653199
transform 1 0 1372 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1711653199
transform 1 0 1268 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1711653199
transform 1 0 1100 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1711653199
transform 1 0 988 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1711653199
transform 1 0 956 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1711653199
transform 1 0 820 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1711653199
transform 1 0 1236 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1711653199
transform 1 0 1124 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1711653199
transform 1 0 732 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1711653199
transform 1 0 700 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1711653199
transform 1 0 548 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1711653199
transform 1 0 436 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1711653199
transform 1 0 396 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1711653199
transform 1 0 316 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1711653199
transform 1 0 396 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1711653199
transform 1 0 276 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1711653199
transform 1 0 252 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1711653199
transform 1 0 188 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1711653199
transform 1 0 396 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1711653199
transform 1 0 252 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_127
timestamp 1711653199
transform 1 0 356 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1711653199
transform 1 0 332 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1711653199
transform 1 0 3396 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1711653199
transform 1 0 3356 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1711653199
transform 1 0 3116 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1711653199
transform 1 0 3076 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_133
timestamp 1711653199
transform 1 0 3332 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1711653199
transform 1 0 3292 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1711653199
transform 1 0 3108 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1711653199
transform 1 0 2980 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1711653199
transform 1 0 2980 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1711653199
transform 1 0 2844 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1711653199
transform 1 0 2724 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1711653199
transform 1 0 2708 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1711653199
transform 1 0 3020 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1711653199
transform 1 0 2996 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_143
timestamp 1711653199
transform 1 0 2980 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1711653199
transform 1 0 2972 0 1 2985
box -2 -2 2 2
use M2_M1  M2_M1_145
timestamp 1711653199
transform 1 0 2772 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1711653199
transform 1 0 2668 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1711653199
transform 1 0 2636 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1711653199
transform 1 0 2316 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1711653199
transform 1 0 1964 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1711653199
transform 1 0 2420 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1711653199
transform 1 0 2364 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1711653199
transform 1 0 2380 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1711653199
transform 1 0 2156 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1711653199
transform 1 0 2268 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1711653199
transform 1 0 2116 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1711653199
transform 1 0 2524 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1711653199
transform 1 0 2308 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1711653199
transform 1 0 2644 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1711653199
transform 1 0 2644 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1711653199
transform 1 0 2636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_161
timestamp 1711653199
transform 1 0 2548 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1711653199
transform 1 0 2116 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1711653199
transform 1 0 1900 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1711653199
transform 1 0 2276 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1711653199
transform 1 0 1860 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1711653199
transform 1 0 1596 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1711653199
transform 1 0 1580 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1711653199
transform 1 0 1708 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1711653199
transform 1 0 1628 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1711653199
transform 1 0 1444 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1711653199
transform 1 0 1404 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1711653199
transform 1 0 1492 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1711653199
transform 1 0 1340 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1711653199
transform 1 0 780 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1711653199
transform 1 0 772 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1711653199
transform 1 0 660 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1711653199
transform 1 0 596 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1711653199
transform 1 0 924 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1711653199
transform 1 0 892 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1711653199
transform 1 0 892 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1711653199
transform 1 0 884 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1711653199
transform 1 0 860 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1711653199
transform 1 0 860 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1711653199
transform 1 0 604 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1711653199
transform 1 0 540 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1711653199
transform 1 0 508 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1711653199
transform 1 0 388 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1711653199
transform 1 0 540 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1711653199
transform 1 0 460 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1711653199
transform 1 0 172 0 1 2385
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1711653199
transform 1 0 172 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1711653199
transform 1 0 116 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1711653199
transform 1 0 116 0 1 2385
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1711653199
transform 1 0 180 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1711653199
transform 1 0 180 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1711653199
transform 1 0 284 0 1 2455
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1711653199
transform 1 0 284 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1711653199
transform 1 0 244 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1711653199
transform 1 0 244 0 1 2455
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1711653199
transform 1 0 388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1711653199
transform 1 0 332 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1711653199
transform 1 0 1124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1711653199
transform 1 0 1084 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1711653199
transform 1 0 1236 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1711653199
transform 1 0 1124 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1711653199
transform 1 0 1436 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1711653199
transform 1 0 1188 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1711653199
transform 1 0 1596 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1711653199
transform 1 0 1276 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1711653199
transform 1 0 1868 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1711653199
transform 1 0 1604 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1711653199
transform 1 0 2012 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1711653199
transform 1 0 1884 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1711653199
transform 1 0 2116 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1711653199
transform 1 0 2076 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1711653199
transform 1 0 2220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1711653199
transform 1 0 2116 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1711653199
transform 1 0 2052 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_219
timestamp 1711653199
transform 1 0 2020 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1711653199
transform 1 0 2452 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1711653199
transform 1 0 2420 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1711653199
transform 1 0 2252 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1711653199
transform 1 0 2220 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1711653199
transform 1 0 2156 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_225
timestamp 1711653199
transform 1 0 2148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1711653199
transform 1 0 2356 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1711653199
transform 1 0 2356 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1711653199
transform 1 0 2796 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1711653199
transform 1 0 2700 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_230
timestamp 1711653199
transform 1 0 2588 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1711653199
transform 1 0 2588 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1711653199
transform 1 0 2004 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_233
timestamp 1711653199
transform 1 0 1956 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1711653199
transform 1 0 1892 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1711653199
transform 1 0 1892 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1711653199
transform 1 0 1652 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1711653199
transform 1 0 1620 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1711653199
transform 1 0 1788 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1711653199
transform 1 0 1660 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1711653199
transform 1 0 1548 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1711653199
transform 1 0 1452 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_242
timestamp 1711653199
transform 1 0 1380 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1711653199
transform 1 0 1380 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1711653199
transform 1 0 900 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1711653199
transform 1 0 852 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1711653199
transform 1 0 668 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1711653199
transform 1 0 660 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1711653199
transform 1 0 1084 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1711653199
transform 1 0 988 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1711653199
transform 1 0 908 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1711653199
transform 1 0 780 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1711653199
transform 1 0 572 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_253
timestamp 1711653199
transform 1 0 508 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1711653199
transform 1 0 460 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1711653199
transform 1 0 452 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1711653199
transform 1 0 500 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1711653199
transform 1 0 364 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1711653199
transform 1 0 172 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1711653199
transform 1 0 172 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_260
timestamp 1711653199
transform 1 0 236 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1711653199
transform 1 0 196 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1711653199
transform 1 0 284 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1711653199
transform 1 0 196 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1711653199
transform 1 0 364 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1711653199
transform 1 0 324 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1711653199
transform 1 0 1116 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1711653199
transform 1 0 508 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1711653199
transform 1 0 1164 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1711653199
transform 1 0 436 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1711653199
transform 1 0 1220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1711653199
transform 1 0 828 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1711653199
transform 1 0 1316 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1711653199
transform 1 0 1076 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1711653199
transform 1 0 1636 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1711653199
transform 1 0 1596 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1711653199
transform 1 0 1916 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1711653199
transform 1 0 1876 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1711653199
transform 1 0 2108 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1711653199
transform 1 0 1940 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_280
timestamp 1711653199
transform 1 0 2148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1711653199
transform 1 0 2068 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1711653199
transform 1 0 3212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1711653199
transform 1 0 3180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1711653199
transform 1 0 3052 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1711653199
transform 1 0 3020 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1711653199
transform 1 0 2924 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1711653199
transform 1 0 2660 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1711653199
transform 1 0 3276 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1711653199
transform 1 0 3252 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1711653199
transform 1 0 3236 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1711653199
transform 1 0 3220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1711653199
transform 1 0 3036 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1711653199
transform 1 0 2996 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1711653199
transform 1 0 2940 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1711653199
transform 1 0 2900 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1711653199
transform 1 0 2516 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1711653199
transform 1 0 2844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1711653199
transform 1 0 2844 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1711653199
transform 1 0 2812 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1711653199
transform 1 0 2500 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1711653199
transform 1 0 2812 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1711653199
transform 1 0 2788 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1711653199
transform 1 0 2772 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1711653199
transform 1 0 2716 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1711653199
transform 1 0 2708 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1711653199
transform 1 0 2548 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1711653199
transform 1 0 2868 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1711653199
transform 1 0 2740 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1711653199
transform 1 0 2700 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1711653199
transform 1 0 2684 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1711653199
transform 1 0 2612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1711653199
transform 1 0 3380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1711653199
transform 1 0 3356 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1711653199
transform 1 0 3316 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1711653199
transform 1 0 3316 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1711653199
transform 1 0 3164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1711653199
transform 1 0 3124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1711653199
transform 1 0 3028 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1711653199
transform 1 0 3316 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1711653199
transform 1 0 3252 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1711653199
transform 1 0 3220 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1711653199
transform 1 0 3212 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_323
timestamp 1711653199
transform 1 0 3204 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1711653199
transform 1 0 3348 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1711653199
transform 1 0 3204 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1711653199
transform 1 0 3196 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_327
timestamp 1711653199
transform 1 0 3188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1711653199
transform 1 0 3068 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1711653199
transform 1 0 3068 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1711653199
transform 1 0 3148 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1711653199
transform 1 0 3020 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1711653199
transform 1 0 3252 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_333
timestamp 1711653199
transform 1 0 3244 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1711653199
transform 1 0 2948 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1711653199
transform 1 0 2820 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1711653199
transform 1 0 2924 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1711653199
transform 1 0 2788 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_338
timestamp 1711653199
transform 1 0 2956 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1711653199
transform 1 0 2844 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1711653199
transform 1 0 3396 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1711653199
transform 1 0 3300 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1711653199
transform 1 0 3260 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1711653199
transform 1 0 3260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1711653199
transform 1 0 3228 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1711653199
transform 1 0 3156 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1711653199
transform 1 0 3140 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1711653199
transform 1 0 3140 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1711653199
transform 1 0 3084 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1711653199
transform 1 0 3036 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1711653199
transform 1 0 3220 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1711653199
transform 1 0 3220 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1711653199
transform 1 0 3196 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1711653199
transform 1 0 3180 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1711653199
transform 1 0 3180 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1711653199
transform 1 0 3140 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1711653199
transform 1 0 3100 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1711653199
transform 1 0 3388 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1711653199
transform 1 0 3252 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1711653199
transform 1 0 3244 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1711653199
transform 1 0 3172 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1711653199
transform 1 0 3172 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1711653199
transform 1 0 3084 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1711653199
transform 1 0 3060 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1711653199
transform 1 0 3052 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1711653199
transform 1 0 2740 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1711653199
transform 1 0 2740 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1711653199
transform 1 0 2964 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1711653199
transform 1 0 2836 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1711653199
transform 1 0 2740 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1711653199
transform 1 0 3052 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1711653199
transform 1 0 2972 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1711653199
transform 1 0 2932 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1711653199
transform 1 0 2932 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1711653199
transform 1 0 3212 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1711653199
transform 1 0 3204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1711653199
transform 1 0 3164 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1711653199
transform 1 0 3164 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1711653199
transform 1 0 3124 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1711653199
transform 1 0 2916 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1711653199
transform 1 0 2916 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1711653199
transform 1 0 2772 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1711653199
transform 1 0 2756 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1711653199
transform 1 0 3236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1711653199
transform 1 0 3180 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1711653199
transform 1 0 3132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1711653199
transform 1 0 3132 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1711653199
transform 1 0 3252 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1711653199
transform 1 0 3252 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1711653199
transform 1 0 3044 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1711653199
transform 1 0 2212 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1711653199
transform 1 0 2108 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1711653199
transform 1 0 2028 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1711653199
transform 1 0 1900 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1711653199
transform 1 0 1660 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1711653199
transform 1 0 1628 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1711653199
transform 1 0 1564 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1711653199
transform 1 0 772 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1711653199
transform 1 0 540 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1711653199
transform 1 0 380 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1711653199
transform 1 0 292 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1711653199
transform 1 0 268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1711653199
transform 1 0 244 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1711653199
transform 1 0 3068 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1711653199
transform 1 0 2836 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1711653199
transform 1 0 2612 0 1 2045
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1711653199
transform 1 0 2580 0 1 2045
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1711653199
transform 1 0 2452 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1711653199
transform 1 0 2364 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1711653199
transform 1 0 2348 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1711653199
transform 1 0 2164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1711653199
transform 1 0 1844 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1711653199
transform 1 0 1844 0 1 2155
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1711653199
transform 1 0 1844 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1711653199
transform 1 0 1828 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1711653199
transform 1 0 1780 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1711653199
transform 1 0 1172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1711653199
transform 1 0 948 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1711653199
transform 1 0 948 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1711653199
transform 1 0 716 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1711653199
transform 1 0 716 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1711653199
transform 1 0 684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1711653199
transform 1 0 660 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_423
timestamp 1711653199
transform 1 0 660 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1711653199
transform 1 0 1532 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1711653199
transform 1 0 1276 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1711653199
transform 1 0 1084 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1711653199
transform 1 0 2892 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1711653199
transform 1 0 2828 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1711653199
transform 1 0 2820 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1711653199
transform 1 0 2788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1711653199
transform 1 0 2748 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1711653199
transform 1 0 2676 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1711653199
transform 1 0 2676 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1711653199
transform 1 0 1716 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1711653199
transform 1 0 1684 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1711653199
transform 1 0 1684 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1711653199
transform 1 0 1652 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1711653199
transform 1 0 1652 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1711653199
transform 1 0 1636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1711653199
transform 1 0 1636 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1711653199
transform 1 0 1572 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1711653199
transform 1 0 1572 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1711653199
transform 1 0 2852 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1711653199
transform 1 0 2772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1711653199
transform 1 0 2684 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1711653199
transform 1 0 2988 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1711653199
transform 1 0 2940 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1711653199
transform 1 0 2836 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1711653199
transform 1 0 2820 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1711653199
transform 1 0 2812 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1711653199
transform 1 0 2804 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1711653199
transform 1 0 2804 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1711653199
transform 1 0 2764 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1711653199
transform 1 0 2748 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1711653199
transform 1 0 2716 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1711653199
transform 1 0 2652 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1711653199
transform 1 0 2308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1711653199
transform 1 0 1332 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1711653199
transform 1 0 1324 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1711653199
transform 1 0 2612 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1711653199
transform 1 0 2612 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1711653199
transform 1 0 2548 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1711653199
transform 1 0 2492 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1711653199
transform 1 0 2436 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1711653199
transform 1 0 2420 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1711653199
transform 1 0 2340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1711653199
transform 1 0 2340 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1711653199
transform 1 0 2332 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1711653199
transform 1 0 2300 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_470
timestamp 1711653199
transform 1 0 2220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1711653199
transform 1 0 2204 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_472
timestamp 1711653199
transform 1 0 2204 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1711653199
transform 1 0 2028 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1711653199
transform 1 0 972 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1711653199
transform 1 0 884 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1711653199
transform 1 0 516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1711653199
transform 1 0 348 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_478
timestamp 1711653199
transform 1 0 332 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1711653199
transform 1 0 212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1711653199
transform 1 0 196 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1711653199
transform 1 0 1788 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1711653199
transform 1 0 1724 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_483
timestamp 1711653199
transform 1 0 1548 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1711653199
transform 1 0 1524 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1711653199
transform 1 0 1476 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1711653199
transform 1 0 1380 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1711653199
transform 1 0 1316 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_488
timestamp 1711653199
transform 1 0 2956 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1711653199
transform 1 0 2932 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1711653199
transform 1 0 2924 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1711653199
transform 1 0 2876 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1711653199
transform 1 0 2868 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1711653199
transform 1 0 2820 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1711653199
transform 1 0 2300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1711653199
transform 1 0 2252 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1711653199
transform 1 0 2252 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1711653199
transform 1 0 2988 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1711653199
transform 1 0 2988 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1711653199
transform 1 0 2948 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1711653199
transform 1 0 2892 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_501
timestamp 1711653199
transform 1 0 2884 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1711653199
transform 1 0 2860 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1711653199
transform 1 0 2860 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1711653199
transform 1 0 2908 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1711653199
transform 1 0 2908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1711653199
transform 1 0 2884 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1711653199
transform 1 0 2852 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1711653199
transform 1 0 2852 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1711653199
transform 1 0 2852 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_510
timestamp 1711653199
transform 1 0 708 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1711653199
transform 1 0 700 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1711653199
transform 1 0 692 0 1 1295
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1711653199
transform 1 0 668 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1711653199
transform 1 0 660 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1711653199
transform 1 0 516 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_516
timestamp 1711653199
transform 1 0 516 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1711653199
transform 1 0 508 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1711653199
transform 1 0 508 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1711653199
transform 1 0 428 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1711653199
transform 1 0 3404 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_521
timestamp 1711653199
transform 1 0 3340 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1711653199
transform 1 0 3044 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1711653199
transform 1 0 3020 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1711653199
transform 1 0 3012 0 1 5
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1711653199
transform 1 0 1468 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1711653199
transform 1 0 1212 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1711653199
transform 1 0 1196 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1711653199
transform 1 0 1172 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1711653199
transform 1 0 1036 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1711653199
transform 1 0 636 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1711653199
transform 1 0 620 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1711653199
transform 1 0 612 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1711653199
transform 1 0 612 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1711653199
transform 1 0 572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1711653199
transform 1 0 548 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1711653199
transform 1 0 484 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1711653199
transform 1 0 92 0 1 85
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1711653199
transform 1 0 3236 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1711653199
transform 1 0 3228 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1711653199
transform 1 0 3180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1711653199
transform 1 0 3140 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1711653199
transform 1 0 2588 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1711653199
transform 1 0 2516 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1711653199
transform 1 0 2516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1711653199
transform 1 0 2468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1711653199
transform 1 0 2452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1711653199
transform 1 0 2356 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1711653199
transform 1 0 2044 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1711653199
transform 1 0 2036 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_550
timestamp 1711653199
transform 1 0 1988 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1711653199
transform 1 0 1988 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1711653199
transform 1 0 1908 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1711653199
transform 1 0 1340 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1711653199
transform 1 0 1324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1711653199
transform 1 0 716 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1711653199
transform 1 0 700 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1711653199
transform 1 0 676 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_558
timestamp 1711653199
transform 1 0 604 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1711653199
transform 1 0 564 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1711653199
transform 1 0 500 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1711653199
transform 1 0 492 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_562
timestamp 1711653199
transform 1 0 1228 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1711653199
transform 1 0 1164 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1711653199
transform 1 0 876 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1711653199
transform 1 0 844 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1711653199
transform 1 0 804 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_567
timestamp 1711653199
transform 1 0 748 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1711653199
transform 1 0 740 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1711653199
transform 1 0 3052 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_570
timestamp 1711653199
transform 1 0 2964 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_571
timestamp 1711653199
transform 1 0 2964 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1711653199
transform 1 0 2956 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1711653199
transform 1 0 2948 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1711653199
transform 1 0 2908 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1711653199
transform 1 0 2908 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1711653199
transform 1 0 1396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1711653199
transform 1 0 2652 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1711653199
transform 1 0 2644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1711653199
transform 1 0 2620 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_580
timestamp 1711653199
transform 1 0 2212 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_581
timestamp 1711653199
transform 1 0 2196 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1711653199
transform 1 0 2180 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1711653199
transform 1 0 2092 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1711653199
transform 1 0 1940 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1711653199
transform 1 0 1836 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1711653199
transform 1 0 2204 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1711653199
transform 1 0 2196 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1711653199
transform 1 0 2172 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1711653199
transform 1 0 2156 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1711653199
transform 1 0 1980 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1711653199
transform 1 0 1980 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1711653199
transform 1 0 1948 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1711653199
transform 1 0 652 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1711653199
transform 1 0 420 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1711653199
transform 1 0 172 0 1 755
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1711653199
transform 1 0 132 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1711653199
transform 1 0 108 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1711653199
transform 1 0 108 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1711653199
transform 1 0 2236 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1711653199
transform 1 0 1844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1711653199
transform 1 0 1812 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1711653199
transform 1 0 1804 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1711653199
transform 1 0 1484 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1711653199
transform 1 0 956 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1711653199
transform 1 0 268 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1711653199
transform 1 0 260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1711653199
transform 1 0 196 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1711653199
transform 1 0 3364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1711653199
transform 1 0 3348 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1711653199
transform 1 0 3332 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1711653199
transform 1 0 3108 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1711653199
transform 1 0 3004 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1711653199
transform 1 0 2940 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1711653199
transform 1 0 2588 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1711653199
transform 1 0 1908 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1711653199
transform 1 0 3116 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1711653199
transform 1 0 2804 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1711653199
transform 1 0 2684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1711653199
transform 1 0 2316 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1711653199
transform 1 0 2300 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1711653199
transform 1 0 2300 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1711653199
transform 1 0 1580 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1711653199
transform 1 0 1092 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1711653199
transform 1 0 1044 0 1 1085
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1711653199
transform 1 0 1028 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1711653199
transform 1 0 1004 0 1 495
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1711653199
transform 1 0 988 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1711653199
transform 1 0 2876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1711653199
transform 1 0 2836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1711653199
transform 1 0 2812 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1711653199
transform 1 0 2788 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1711653199
transform 1 0 2764 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1711653199
transform 1 0 2636 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1711653199
transform 1 0 2636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1711653199
transform 1 0 2580 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1711653199
transform 1 0 2524 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1711653199
transform 1 0 2020 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1711653199
transform 1 0 2020 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1711653199
transform 1 0 2620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1711653199
transform 1 0 2596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1711653199
transform 1 0 2588 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1711653199
transform 1 0 2556 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1711653199
transform 1 0 2556 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1711653199
transform 1 0 2540 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1711653199
transform 1 0 2260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1711653199
transform 1 0 2228 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1711653199
transform 1 0 2228 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1711653199
transform 1 0 348 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1711653199
transform 1 0 300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1711653199
transform 1 0 2140 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1711653199
transform 1 0 2140 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1711653199
transform 1 0 2108 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1711653199
transform 1 0 2100 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1711653199
transform 1 0 2084 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1711653199
transform 1 0 2076 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1711653199
transform 1 0 1900 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1711653199
transform 1 0 1628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1711653199
transform 1 0 1604 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1711653199
transform 1 0 1076 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1711653199
transform 1 0 500 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1711653199
transform 1 0 436 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1711653199
transform 1 0 2756 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1711653199
transform 1 0 2724 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1711653199
transform 1 0 2676 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1711653199
transform 1 0 2612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1711653199
transform 1 0 2540 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1711653199
transform 1 0 2276 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1711653199
transform 1 0 2276 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1711653199
transform 1 0 2252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1711653199
transform 1 0 2252 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1711653199
transform 1 0 2228 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1711653199
transform 1 0 1548 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1711653199
transform 1 0 2612 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1711653199
transform 1 0 2612 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1711653199
transform 1 0 2556 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1711653199
transform 1 0 2532 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1711653199
transform 1 0 1012 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1711653199
transform 1 0 1004 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1711653199
transform 1 0 940 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1711653199
transform 1 0 932 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1711653199
transform 1 0 860 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1711653199
transform 1 0 2668 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1711653199
transform 1 0 2660 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1711653199
transform 1 0 2308 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1711653199
transform 1 0 2292 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1711653199
transform 1 0 2044 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1711653199
transform 1 0 2004 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1711653199
transform 1 0 1372 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1711653199
transform 1 0 1204 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1711653199
transform 1 0 1204 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1711653199
transform 1 0 1196 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1711653199
transform 1 0 1196 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1711653199
transform 1 0 1164 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1711653199
transform 1 0 1148 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1711653199
transform 1 0 436 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1711653199
transform 1 0 404 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1711653199
transform 1 0 396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1711653199
transform 1 0 388 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1711653199
transform 1 0 380 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1711653199
transform 1 0 340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1711653199
transform 1 0 580 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1711653199
transform 1 0 564 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1711653199
transform 1 0 516 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1711653199
transform 1 0 484 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1711653199
transform 1 0 444 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1711653199
transform 1 0 348 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_707
timestamp 1711653199
transform 1 0 252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1711653199
transform 1 0 228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1711653199
transform 1 0 148 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1711653199
transform 1 0 108 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1711653199
transform 1 0 3372 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1711653199
transform 1 0 3364 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1711653199
transform 1 0 3356 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1711653199
transform 1 0 3332 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1711653199
transform 1 0 3316 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1711653199
transform 1 0 1372 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1711653199
transform 1 0 1364 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1711653199
transform 1 0 1300 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1711653199
transform 1 0 1276 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1711653199
transform 1 0 1252 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1711653199
transform 1 0 1204 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1711653199
transform 1 0 1140 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1711653199
transform 1 0 1132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1711653199
transform 1 0 3196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1711653199
transform 1 0 3196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1711653199
transform 1 0 3108 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1711653199
transform 1 0 3092 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1711653199
transform 1 0 3052 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1711653199
transform 1 0 2612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1711653199
transform 1 0 2556 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1711653199
transform 1 0 2556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1711653199
transform 1 0 2532 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1711653199
transform 1 0 2524 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1711653199
transform 1 0 2300 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1711653199
transform 1 0 2300 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_736
timestamp 1711653199
transform 1 0 2284 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_737
timestamp 1711653199
transform 1 0 3316 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_738
timestamp 1711653199
transform 1 0 3308 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1711653199
transform 1 0 3308 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1711653199
transform 1 0 3284 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_741
timestamp 1711653199
transform 1 0 3268 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1711653199
transform 1 0 2412 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1711653199
transform 1 0 2212 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1711653199
transform 1 0 372 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1711653199
transform 1 0 364 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_746
timestamp 1711653199
transform 1 0 348 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1711653199
transform 1 0 332 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1711653199
transform 1 0 324 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1711653199
transform 1 0 316 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1711653199
transform 1 0 316 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1711653199
transform 1 0 316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1711653199
transform 1 0 308 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1711653199
transform 1 0 308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1711653199
transform 1 0 284 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1711653199
transform 1 0 276 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1711653199
transform 1 0 220 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_757
timestamp 1711653199
transform 1 0 212 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1711653199
transform 1 0 3380 0 1 1185
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1711653199
transform 1 0 3300 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1711653199
transform 1 0 3292 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1711653199
transform 1 0 3220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1711653199
transform 1 0 3220 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1711653199
transform 1 0 3180 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1711653199
transform 1 0 2604 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1711653199
transform 1 0 2148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_766
timestamp 1711653199
transform 1 0 356 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1711653199
transform 1 0 340 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1711653199
transform 1 0 300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1711653199
transform 1 0 300 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1711653199
transform 1 0 300 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1711653199
transform 1 0 292 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_772
timestamp 1711653199
transform 1 0 292 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1711653199
transform 1 0 276 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1711653199
transform 1 0 260 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1711653199
transform 1 0 236 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1711653199
transform 1 0 196 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1711653199
transform 1 0 2180 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1711653199
transform 1 0 2164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1711653199
transform 1 0 2044 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1711653199
transform 1 0 1852 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1711653199
transform 1 0 1836 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1711653199
transform 1 0 1412 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1711653199
transform 1 0 1372 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1711653199
transform 1 0 1324 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1711653199
transform 1 0 628 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1711653199
transform 1 0 428 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1711653199
transform 1 0 308 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1711653199
transform 1 0 268 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1711653199
transform 1 0 268 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1711653199
transform 1 0 236 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_791
timestamp 1711653199
transform 1 0 236 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1711653199
transform 1 0 196 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1711653199
transform 1 0 1164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1711653199
transform 1 0 1084 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1711653199
transform 1 0 1020 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1711653199
transform 1 0 820 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1711653199
transform 1 0 620 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1711653199
transform 1 0 452 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1711653199
transform 1 0 436 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1711653199
transform 1 0 404 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1711653199
transform 1 0 396 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1711653199
transform 1 0 3364 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1711653199
transform 1 0 3356 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1711653199
transform 1 0 3356 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1711653199
transform 1 0 3252 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1711653199
transform 1 0 2860 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1711653199
transform 1 0 2860 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1711653199
transform 1 0 2772 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_809
timestamp 1711653199
transform 1 0 1348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1711653199
transform 1 0 2612 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1711653199
transform 1 0 2596 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1711653199
transform 1 0 2580 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1711653199
transform 1 0 2244 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1711653199
transform 1 0 2092 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1711653199
transform 1 0 2028 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1711653199
transform 1 0 1708 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1711653199
transform 1 0 1260 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1711653199
transform 1 0 1252 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1711653199
transform 1 0 1252 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1711653199
transform 1 0 1220 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1711653199
transform 1 0 1156 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1711653199
transform 1 0 532 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1711653199
transform 1 0 484 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1711653199
transform 1 0 420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1711653199
transform 1 0 412 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1711653199
transform 1 0 388 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1711653199
transform 1 0 2220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1711653199
transform 1 0 2204 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1711653199
transform 1 0 2092 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1711653199
transform 1 0 1948 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1711653199
transform 1 0 1620 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_832
timestamp 1711653199
transform 1 0 1492 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1711653199
transform 1 0 1484 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1711653199
transform 1 0 1476 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1711653199
transform 1 0 788 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1711653199
transform 1 0 708 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1711653199
transform 1 0 2908 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1711653199
transform 1 0 2556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1711653199
transform 1 0 2516 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1711653199
transform 1 0 2492 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1711653199
transform 1 0 2292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1711653199
transform 1 0 1916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1711653199
transform 1 0 2972 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1711653199
transform 1 0 2868 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1711653199
transform 1 0 2316 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1711653199
transform 1 0 1388 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1711653199
transform 1 0 1380 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1711653199
transform 1 0 1300 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1711653199
transform 1 0 1204 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1711653199
transform 1 0 1164 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1711653199
transform 1 0 1108 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1711653199
transform 1 0 1060 0 1 1185
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1711653199
transform 1 0 1020 0 1 1245
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1711653199
transform 1 0 1020 0 1 1185
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1711653199
transform 1 0 972 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1711653199
transform 1 0 972 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1711653199
transform 1 0 948 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1711653199
transform 1 0 2564 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1711653199
transform 1 0 2508 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1711653199
transform 1 0 2436 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1711653199
transform 1 0 2436 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1711653199
transform 1 0 2876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1711653199
transform 1 0 2788 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1711653199
transform 1 0 2772 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1711653199
transform 1 0 2668 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_866
timestamp 1711653199
transform 1 0 2452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1711653199
transform 1 0 2452 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1711653199
transform 1 0 2436 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1711653199
transform 1 0 2436 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1711653199
transform 1 0 2436 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1711653199
transform 1 0 2396 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1711653199
transform 1 0 2372 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1711653199
transform 1 0 1860 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1711653199
transform 1 0 1860 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1711653199
transform 1 0 1860 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1711653199
transform 1 0 1676 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1711653199
transform 1 0 884 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1711653199
transform 1 0 868 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1711653199
transform 1 0 2332 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1711653199
transform 1 0 2324 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1711653199
transform 1 0 2276 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1711653199
transform 1 0 1932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1711653199
transform 1 0 1916 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1711653199
transform 1 0 3060 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1711653199
transform 1 0 3060 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1711653199
transform 1 0 2444 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1711653199
transform 1 0 2100 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1711653199
transform 1 0 1836 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1711653199
transform 1 0 1012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1711653199
transform 1 0 980 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1711653199
transform 1 0 964 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1711653199
transform 1 0 908 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1711653199
transform 1 0 892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1711653199
transform 1 0 764 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1711653199
transform 1 0 716 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1711653199
transform 1 0 636 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1711653199
transform 1 0 628 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1711653199
transform 1 0 2140 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1711653199
transform 1 0 2100 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1711653199
transform 1 0 2084 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1711653199
transform 1 0 2460 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1711653199
transform 1 0 2460 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1711653199
transform 1 0 2444 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1711653199
transform 1 0 2420 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1711653199
transform 1 0 2420 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1711653199
transform 1 0 2388 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1711653199
transform 1 0 2388 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1711653199
transform 1 0 2364 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1711653199
transform 1 0 2364 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1711653199
transform 1 0 2340 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1711653199
transform 1 0 2332 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1711653199
transform 1 0 2324 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1711653199
transform 1 0 2308 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1711653199
transform 1 0 2308 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1711653199
transform 1 0 1652 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1711653199
transform 1 0 1548 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1711653199
transform 1 0 1476 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1711653199
transform 1 0 1244 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1711653199
transform 1 0 1220 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1711653199
transform 1 0 1220 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1711653199
transform 1 0 1196 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1711653199
transform 1 0 980 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1711653199
transform 1 0 892 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1711653199
transform 1 0 884 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_925
timestamp 1711653199
transform 1 0 884 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1711653199
transform 1 0 868 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1711653199
transform 1 0 868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_928
timestamp 1711653199
transform 1 0 852 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1711653199
transform 1 0 852 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1711653199
transform 1 0 796 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1711653199
transform 1 0 788 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1711653199
transform 1 0 692 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1711653199
transform 1 0 612 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1711653199
transform 1 0 2100 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1711653199
transform 1 0 2100 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1711653199
transform 1 0 2060 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1711653199
transform 1 0 2140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1711653199
transform 1 0 2116 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_939
timestamp 1711653199
transform 1 0 2076 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1711653199
transform 1 0 1988 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1711653199
transform 1 0 1860 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1711653199
transform 1 0 1708 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1711653199
transform 1 0 1660 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1711653199
transform 1 0 1644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1711653199
transform 1 0 1628 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1711653199
transform 1 0 1564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1711653199
transform 1 0 1556 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1711653199
transform 1 0 1556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1711653199
transform 1 0 1556 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1711653199
transform 1 0 1548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1711653199
transform 1 0 1548 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1711653199
transform 1 0 1516 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1711653199
transform 1 0 1508 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1711653199
transform 1 0 1340 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1711653199
transform 1 0 1292 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1711653199
transform 1 0 1260 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1711653199
transform 1 0 2308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1711653199
transform 1 0 2212 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1711653199
transform 1 0 2196 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1711653199
transform 1 0 2172 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1711653199
transform 1 0 2108 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1711653199
transform 1 0 1636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1711653199
transform 1 0 1532 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1711653199
transform 1 0 1252 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1711653199
transform 1 0 1220 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1711653199
transform 1 0 1180 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1711653199
transform 1 0 1132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1711653199
transform 1 0 1084 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1711653199
transform 1 0 1068 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1711653199
transform 1 0 1060 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1711653199
transform 1 0 940 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1711653199
transform 1 0 916 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1711653199
transform 1 0 868 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1711653199
transform 1 0 2396 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1711653199
transform 1 0 2364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1711653199
transform 1 0 2268 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1711653199
transform 1 0 2268 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1711653199
transform 1 0 2212 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1711653199
transform 1 0 2204 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1711653199
transform 1 0 2436 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1711653199
transform 1 0 2356 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_982
timestamp 1711653199
transform 1 0 2356 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1711653199
transform 1 0 2340 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1711653199
transform 1 0 2236 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1711653199
transform 1 0 2196 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1711653199
transform 1 0 1908 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1711653199
transform 1 0 1900 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1711653199
transform 1 0 1028 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1711653199
transform 1 0 916 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1711653199
transform 1 0 876 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1711653199
transform 1 0 860 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1711653199
transform 1 0 812 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1711653199
transform 1 0 780 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1711653199
transform 1 0 500 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1711653199
transform 1 0 3068 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1711653199
transform 1 0 2332 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1711653199
transform 1 0 1540 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1711653199
transform 1 0 1492 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1711653199
transform 1 0 1364 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1711653199
transform 1 0 1188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1001
timestamp 1711653199
transform 1 0 700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1711653199
transform 1 0 508 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1711653199
transform 1 0 444 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1711653199
transform 1 0 404 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1711653199
transform 1 0 380 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1711653199
transform 1 0 3292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1007
timestamp 1711653199
transform 1 0 3268 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1711653199
transform 1 0 3204 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1711653199
transform 1 0 3148 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1711653199
transform 1 0 2972 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1011
timestamp 1711653199
transform 1 0 2916 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1711653199
transform 1 0 2708 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1711653199
transform 1 0 2636 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1711653199
transform 1 0 2620 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1015
timestamp 1711653199
transform 1 0 2612 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1711653199
transform 1 0 1772 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1711653199
transform 1 0 1756 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1711653199
transform 1 0 1252 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1711653199
transform 1 0 1188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1711653199
transform 1 0 1124 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1711653199
transform 1 0 588 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1711653199
transform 1 0 292 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1023
timestamp 1711653199
transform 1 0 236 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1711653199
transform 1 0 220 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1711653199
transform 1 0 204 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1711653199
transform 1 0 164 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1711653199
transform 1 0 476 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1711653199
transform 1 0 452 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1711653199
transform 1 0 420 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1711653199
transform 1 0 340 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1711653199
transform 1 0 3396 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1711653199
transform 1 0 3340 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1711653199
transform 1 0 3212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1711653199
transform 1 0 2732 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1711653199
transform 1 0 2508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1711653199
transform 1 0 2516 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1711653199
transform 1 0 2404 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1711653199
transform 1 0 1732 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1711653199
transform 1 0 1724 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1711653199
transform 1 0 1668 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1711653199
transform 1 0 1660 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1711653199
transform 1 0 1140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1711653199
transform 1 0 1036 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1711653199
transform 1 0 988 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1711653199
transform 1 0 508 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1711653199
transform 1 0 1332 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1711653199
transform 1 0 1260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1711653199
transform 1 0 1236 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1711653199
transform 1 0 2404 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1711653199
transform 1 0 2172 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1711653199
transform 1 0 2084 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1711653199
transform 1 0 2764 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1711653199
transform 1 0 2628 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1711653199
transform 1 0 2532 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1055
timestamp 1711653199
transform 1 0 2524 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1711653199
transform 1 0 1884 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1711653199
transform 1 0 1860 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1711653199
transform 1 0 1836 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1711653199
transform 1 0 1820 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1711653199
transform 1 0 1796 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1711653199
transform 1 0 1756 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1711653199
transform 1 0 1748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1711653199
transform 1 0 2308 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1711653199
transform 1 0 2308 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1711653199
transform 1 0 2260 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1711653199
transform 1 0 2236 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1711653199
transform 1 0 2212 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1711653199
transform 1 0 684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1711653199
transform 1 0 652 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1711653199
transform 1 0 572 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1711653199
transform 1 0 364 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1711653199
transform 1 0 756 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1711653199
transform 1 0 740 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1074
timestamp 1711653199
transform 1 0 676 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1711653199
transform 1 0 540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1711653199
transform 1 0 3276 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1711653199
transform 1 0 3228 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1711653199
transform 1 0 3020 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1711653199
transform 1 0 3012 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1711653199
transform 1 0 1780 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1711653199
transform 1 0 1732 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1711653199
transform 1 0 1692 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1711653199
transform 1 0 1796 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1711653199
transform 1 0 1764 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1711653199
transform 1 0 644 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1711653199
transform 1 0 644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1711653199
transform 1 0 636 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1088
timestamp 1711653199
transform 1 0 596 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1089
timestamp 1711653199
transform 1 0 596 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1711653199
transform 1 0 580 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1711653199
transform 1 0 572 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1711653199
transform 1 0 892 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1711653199
transform 1 0 812 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1711653199
transform 1 0 764 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1711653199
transform 1 0 748 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1711653199
transform 1 0 732 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1711653199
transform 1 0 732 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1711653199
transform 1 0 2540 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1711653199
transform 1 0 2260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1711653199
transform 1 0 1956 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1711653199
transform 1 0 3172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1711653199
transform 1 0 3100 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1103
timestamp 1711653199
transform 1 0 3092 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1711653199
transform 1 0 3004 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1711653199
transform 1 0 2956 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1711653199
transform 1 0 2660 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1711653199
transform 1 0 2628 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1711653199
transform 1 0 2628 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1711653199
transform 1 0 1900 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1711653199
transform 1 0 1892 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1711653199
transform 1 0 1884 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1112
timestamp 1711653199
transform 1 0 1708 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1711653199
transform 1 0 1692 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1711653199
transform 1 0 1684 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1711653199
transform 1 0 2124 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1711653199
transform 1 0 1956 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1711653199
transform 1 0 1956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1711653199
transform 1 0 892 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1711653199
transform 1 0 796 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1711653199
transform 1 0 372 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1711653199
transform 1 0 356 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1711653199
transform 1 0 164 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1711653199
transform 1 0 156 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1124
timestamp 1711653199
transform 1 0 124 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1711653199
transform 1 0 116 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1711653199
transform 1 0 1604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1127
timestamp 1711653199
transform 1 0 1532 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1711653199
transform 1 0 1508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1711653199
transform 1 0 1124 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1711653199
transform 1 0 340 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1711653199
transform 1 0 316 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1132
timestamp 1711653199
transform 1 0 316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1711653199
transform 1 0 268 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1711653199
transform 1 0 3348 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1711653199
transform 1 0 3300 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1711653199
transform 1 0 3300 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1711653199
transform 1 0 3108 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1711653199
transform 1 0 2932 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1711653199
transform 1 0 2908 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1711653199
transform 1 0 2908 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1711653199
transform 1 0 1900 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1711653199
transform 1 0 1860 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1711653199
transform 1 0 1020 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1711653199
transform 1 0 804 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1711653199
transform 1 0 524 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1711653199
transform 1 0 156 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1711653199
transform 1 0 148 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1711653199
transform 1 0 1316 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1711653199
transform 1 0 1236 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1711653199
transform 1 0 636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1711653199
transform 1 0 588 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1711653199
transform 1 0 332 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1711653199
transform 1 0 276 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1711653199
transform 1 0 3396 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1711653199
transform 1 0 3308 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1156
timestamp 1711653199
transform 1 0 2860 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1711653199
transform 1 0 2780 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1711653199
transform 1 0 2476 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1711653199
transform 1 0 2180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1711653199
transform 1 0 1228 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1711653199
transform 1 0 1212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1711653199
transform 1 0 2028 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1711653199
transform 1 0 2004 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1164
timestamp 1711653199
transform 1 0 1844 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1711653199
transform 1 0 1820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1711653199
transform 1 0 1820 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1711653199
transform 1 0 1756 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1711653199
transform 1 0 1796 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1711653199
transform 1 0 1620 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1711653199
transform 1 0 1572 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1711653199
transform 1 0 1508 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1711653199
transform 1 0 1396 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1711653199
transform 1 0 956 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1711653199
transform 1 0 916 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1711653199
transform 1 0 708 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1711653199
transform 1 0 700 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1711653199
transform 1 0 372 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1711653199
transform 1 0 364 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1711653199
transform 1 0 348 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1711653199
transform 1 0 540 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1711653199
transform 1 0 540 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1711653199
transform 1 0 212 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1711653199
transform 1 0 204 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1711653199
transform 1 0 220 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1711653199
transform 1 0 220 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1711653199
transform 1 0 404 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1711653199
transform 1 0 260 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1711653199
transform 1 0 260 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1711653199
transform 1 0 228 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1711653199
transform 1 0 212 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1711653199
transform 1 0 260 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1711653199
transform 1 0 260 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1711653199
transform 1 0 260 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1711653199
transform 1 0 476 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1711653199
transform 1 0 412 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1711653199
transform 1 0 412 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1711653199
transform 1 0 780 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1711653199
transform 1 0 764 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1711653199
transform 1 0 724 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1200
timestamp 1711653199
transform 1 0 708 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1711653199
transform 1 0 1132 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1711653199
transform 1 0 1132 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1711653199
transform 1 0 908 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1711653199
transform 1 0 804 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1711653199
transform 1 0 804 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1711653199
transform 1 0 1012 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1711653199
transform 1 0 972 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1208
timestamp 1711653199
transform 1 0 972 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1711653199
transform 1 0 1300 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1711653199
transform 1 0 1260 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1711653199
transform 1 0 1516 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1711653199
transform 1 0 1492 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1711653199
transform 1 0 1476 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1711653199
transform 1 0 1748 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1711653199
transform 1 0 1708 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1711653199
transform 1 0 1636 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1711653199
transform 1 0 1636 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1711653199
transform 1 0 1596 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1711653199
transform 1 0 1876 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1711653199
transform 1 0 1876 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1221
timestamp 1711653199
transform 1 0 1828 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1711653199
transform 1 0 1948 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1711653199
transform 1 0 1932 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1711653199
transform 1 0 2308 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1711653199
transform 1 0 2276 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1711653199
transform 1 0 2220 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1227
timestamp 1711653199
transform 1 0 2188 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1711653199
transform 1 0 2172 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1711653199
transform 1 0 2492 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1711653199
transform 1 0 2476 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1711653199
transform 1 0 2324 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1711653199
transform 1 0 2436 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1711653199
transform 1 0 2428 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1711653199
transform 1 0 2388 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1711653199
transform 1 0 2044 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1711653199
transform 1 0 2004 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1711653199
transform 1 0 3172 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1711653199
transform 1 0 3156 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1239
timestamp 1711653199
transform 1 0 3116 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1711653199
transform 1 0 2684 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1711653199
transform 1 0 2452 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1711653199
transform 1 0 3292 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1711653199
transform 1 0 3276 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1244
timestamp 1711653199
transform 1 0 3268 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1711653199
transform 1 0 3116 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1711653199
transform 1 0 3116 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1711653199
transform 1 0 3084 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1711653199
transform 1 0 3044 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1711653199
transform 1 0 3044 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1711653199
transform 1 0 3012 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1711653199
transform 1 0 3284 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1711653199
transform 1 0 3140 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1711653199
transform 1 0 3108 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1711653199
transform 1 0 3364 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1711653199
transform 1 0 3252 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1711653199
transform 1 0 3132 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1711653199
transform 1 0 3100 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1711653199
transform 1 0 3364 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1259
timestamp 1711653199
transform 1 0 3252 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1711653199
transform 1 0 3364 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1711653199
transform 1 0 3332 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1711653199
transform 1 0 3228 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1711653199
transform 1 0 3140 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_1264
timestamp 1711653199
transform 1 0 3140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1711653199
transform 1 0 2804 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1711653199
transform 1 0 2788 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1711653199
transform 1 0 2732 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1711653199
transform 1 0 2716 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1711653199
transform 1 0 2780 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1711653199
transform 1 0 2764 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1711653199
transform 1 0 2748 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1711653199
transform 1 0 2988 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1711653199
transform 1 0 2932 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1711653199
transform 1 0 2924 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1711653199
transform 1 0 2916 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1711653199
transform 1 0 2876 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1711653199
transform 1 0 3220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1711653199
transform 1 0 3204 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1711653199
transform 1 0 3180 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1711653199
transform 1 0 3148 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1711653199
transform 1 0 3148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1711653199
transform 1 0 3116 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1711653199
transform 1 0 3116 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1711653199
transform 1 0 3252 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1711653199
transform 1 0 3236 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1711653199
transform 1 0 3204 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1711653199
transform 1 0 3180 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1711653199
transform 1 0 3252 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1711653199
transform 1 0 3228 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1290
timestamp 1711653199
transform 1 0 3220 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1711653199
transform 1 0 3180 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1711653199
transform 1 0 3156 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1711653199
transform 1 0 3140 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1294
timestamp 1711653199
transform 1 0 3132 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1711653199
transform 1 0 3116 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1711653199
transform 1 0 3028 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1711653199
transform 1 0 2964 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1711653199
transform 1 0 2412 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1711653199
transform 1 0 2388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1711653199
transform 1 0 2188 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1711653199
transform 1 0 3228 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1711653199
transform 1 0 3228 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1711653199
transform 1 0 3084 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1711653199
transform 1 0 3044 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1711653199
transform 1 0 1140 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1711653199
transform 1 0 1084 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1711653199
transform 1 0 1068 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1711653199
transform 1 0 972 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1711653199
transform 1 0 964 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1711653199
transform 1 0 980 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1711653199
transform 1 0 964 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1711653199
transform 1 0 2156 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1711653199
transform 1 0 2116 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1711653199
transform 1 0 2412 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1711653199
transform 1 0 2324 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1711653199
transform 1 0 2516 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1711653199
transform 1 0 2500 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1318
timestamp 1711653199
transform 1 0 3036 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1711653199
transform 1 0 2940 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1711653199
transform 1 0 2932 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1711653199
transform 1 0 2988 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1711653199
transform 1 0 2956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1711653199
transform 1 0 3100 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1711653199
transform 1 0 3100 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1711653199
transform 1 0 2996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1711653199
transform 1 0 2996 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1711653199
transform 1 0 2980 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1711653199
transform 1 0 2972 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1711653199
transform 1 0 2956 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1711653199
transform 1 0 3364 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1711653199
transform 1 0 3324 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1711653199
transform 1 0 3324 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1333
timestamp 1711653199
transform 1 0 3340 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_1334
timestamp 1711653199
transform 1 0 3316 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1711653199
transform 1 0 3316 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1711653199
transform 1 0 3356 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1711653199
transform 1 0 3356 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1711653199
transform 1 0 3332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1711653199
transform 1 0 3340 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1711653199
transform 1 0 3116 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1341
timestamp 1711653199
transform 1 0 3396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1711653199
transform 1 0 3324 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1711653199
transform 1 0 3260 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1711653199
transform 1 0 3196 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1711653199
transform 1 0 3172 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1346
timestamp 1711653199
transform 1 0 1468 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1711653199
transform 1 0 1468 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1711653199
transform 1 0 1428 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1711653199
transform 1 0 1372 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1711653199
transform 1 0 2756 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1711653199
transform 1 0 2692 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1711653199
transform 1 0 2668 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1711653199
transform 1 0 2636 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1354
timestamp 1711653199
transform 1 0 2636 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1711653199
transform 1 0 2652 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1711653199
transform 1 0 2628 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1711653199
transform 1 0 2844 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1711653199
transform 1 0 2804 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1711653199
transform 1 0 2716 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1711653199
transform 1 0 2708 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1711653199
transform 1 0 2660 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1711653199
transform 1 0 2636 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1711653199
transform 1 0 2724 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1711653199
transform 1 0 2676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1711653199
transform 1 0 2012 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1711653199
transform 1 0 2124 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1711653199
transform 1 0 2124 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1711653199
transform 1 0 2100 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1711653199
transform 1 0 1956 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1711653199
transform 1 0 1956 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1371
timestamp 1711653199
transform 1 0 1444 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1711653199
transform 1 0 2148 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1711653199
transform 1 0 2148 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1711653199
transform 1 0 1740 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1711653199
transform 1 0 1484 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1711653199
transform 1 0 2332 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1711653199
transform 1 0 2308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1711653199
transform 1 0 2212 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1711653199
transform 1 0 2204 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1711653199
transform 1 0 2060 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1711653199
transform 1 0 2052 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1711653199
transform 1 0 2516 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1711653199
transform 1 0 2468 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1384
timestamp 1711653199
transform 1 0 2372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1385
timestamp 1711653199
transform 1 0 2340 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1711653199
transform 1 0 2364 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1387
timestamp 1711653199
transform 1 0 2292 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1711653199
transform 1 0 2252 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1711653199
transform 1 0 2228 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1711653199
transform 1 0 2604 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1711653199
transform 1 0 2564 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1711653199
transform 1 0 2300 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1393
timestamp 1711653199
transform 1 0 2284 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1711653199
transform 1 0 1220 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1395
timestamp 1711653199
transform 1 0 1220 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1396
timestamp 1711653199
transform 1 0 2276 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1711653199
transform 1 0 2020 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1711653199
transform 1 0 1980 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1711653199
transform 1 0 2364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1400
timestamp 1711653199
transform 1 0 2324 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1711653199
transform 1 0 2540 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_1402
timestamp 1711653199
transform 1 0 2380 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1711653199
transform 1 0 2380 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1711653199
transform 1 0 2564 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1711653199
transform 1 0 2564 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1711653199
transform 1 0 2148 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1711653199
transform 1 0 2140 0 1 1495
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1711653199
transform 1 0 2076 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1711653199
transform 1 0 2060 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1410
timestamp 1711653199
transform 1 0 2060 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1711653199
transform 1 0 2156 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1711653199
transform 1 0 2084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1711653199
transform 1 0 2084 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1711653199
transform 1 0 1764 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1711653199
transform 1 0 1748 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1711653199
transform 1 0 1788 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1417
timestamp 1711653199
transform 1 0 1788 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1711653199
transform 1 0 2508 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1711653199
transform 1 0 1940 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1711653199
transform 1 0 1940 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1421
timestamp 1711653199
transform 1 0 1684 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1711653199
transform 1 0 1532 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1711653199
transform 1 0 1292 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1424
timestamp 1711653199
transform 1 0 1868 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1711653199
transform 1 0 1868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1426
timestamp 1711653199
transform 1 0 2228 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1711653199
transform 1 0 1820 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1428
timestamp 1711653199
transform 1 0 1796 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1711653199
transform 1 0 1508 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1430
timestamp 1711653199
transform 1 0 1508 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1711653199
transform 1 0 1468 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1711653199
transform 1 0 1468 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_1433
timestamp 1711653199
transform 1 0 1428 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1711653199
transform 1 0 1428 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1711653199
transform 1 0 1148 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1711653199
transform 1 0 1060 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1711653199
transform 1 0 1036 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1711653199
transform 1 0 2036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1711653199
transform 1 0 2004 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1711653199
transform 1 0 2188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1711653199
transform 1 0 2172 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1711653199
transform 1 0 756 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1711653199
transform 1 0 756 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1711653199
transform 1 0 684 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1711653199
transform 1 0 644 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1711653199
transform 1 0 604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1711653199
transform 1 0 772 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1711653199
transform 1 0 700 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1711653199
transform 1 0 700 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1711653199
transform 1 0 628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1711653199
transform 1 0 612 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1711653199
transform 1 0 260 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1711653199
transform 1 0 252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1711653199
transform 1 0 228 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1711653199
transform 1 0 332 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1711653199
transform 1 0 260 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_1457
timestamp 1711653199
transform 1 0 228 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1711653199
transform 1 0 196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1711653199
transform 1 0 188 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_1460
timestamp 1711653199
transform 1 0 180 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1711653199
transform 1 0 164 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1711653199
transform 1 0 164 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1711653199
transform 1 0 116 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1464
timestamp 1711653199
transform 1 0 108 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1711653199
transform 1 0 92 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1711653199
transform 1 0 84 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1711653199
transform 1 0 180 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1711653199
transform 1 0 132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1711653199
transform 1 0 100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1711653199
transform 1 0 100 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_1471
timestamp 1711653199
transform 1 0 92 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1711653199
transform 1 0 68 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1473
timestamp 1711653199
transform 1 0 68 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1711653199
transform 1 0 1204 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1711653199
transform 1 0 1180 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1711653199
transform 1 0 1156 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_1477
timestamp 1711653199
transform 1 0 1140 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1711653199
transform 1 0 1092 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1711653199
transform 1 0 1068 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1711653199
transform 1 0 868 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1711653199
transform 1 0 860 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1711653199
transform 1 0 708 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1711653199
transform 1 0 676 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1711653199
transform 1 0 644 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1711653199
transform 1 0 996 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1711653199
transform 1 0 948 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1711653199
transform 1 0 916 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1711653199
transform 1 0 1260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1489
timestamp 1711653199
transform 1 0 1220 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1711653199
transform 1 0 972 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1711653199
transform 1 0 468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1711653199
transform 1 0 468 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1711653199
transform 1 0 948 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1711653199
transform 1 0 892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1711653199
transform 1 0 828 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1711653199
transform 1 0 700 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_1497
timestamp 1711653199
transform 1 0 860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1711653199
transform 1 0 812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1711653199
transform 1 0 692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1711653199
transform 1 0 676 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1711653199
transform 1 0 652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1711653199
transform 1 0 588 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1711653199
transform 1 0 1260 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_1504
timestamp 1711653199
transform 1 0 644 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1711653199
transform 1 0 580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1711653199
transform 1 0 492 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1507
timestamp 1711653199
transform 1 0 436 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1508
timestamp 1711653199
transform 1 0 1116 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1711653199
transform 1 0 860 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1711653199
transform 1 0 596 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1711653199
transform 1 0 996 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1512
timestamp 1711653199
transform 1 0 756 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1711653199
transform 1 0 596 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1711653199
transform 1 0 572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1711653199
transform 1 0 1124 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1711653199
transform 1 0 1124 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1711653199
transform 1 0 1092 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1711653199
transform 1 0 956 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1519
timestamp 1711653199
transform 1 0 932 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1711653199
transform 1 0 2372 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1711653199
transform 1 0 2372 0 1 555
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1711653199
transform 1 0 1772 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1711653199
transform 1 0 1772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1711653199
transform 1 0 852 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1711653199
transform 1 0 844 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1711653199
transform 1 0 1052 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1711653199
transform 1 0 996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1711653199
transform 1 0 1052 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1711653199
transform 1 0 900 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1711653199
transform 1 0 900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1531
timestamp 1711653199
transform 1 0 964 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1711653199
transform 1 0 892 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1533
timestamp 1711653199
transform 1 0 772 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1711653199
transform 1 0 756 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1711653199
transform 1 0 452 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1711653199
transform 1 0 452 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1711653199
transform 1 0 436 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1538
timestamp 1711653199
transform 1 0 428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1711653199
transform 1 0 428 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1711653199
transform 1 0 412 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1711653199
transform 1 0 364 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1711653199
transform 1 0 364 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1711653199
transform 1 0 124 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1711653199
transform 1 0 76 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1711653199
transform 1 0 228 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1711653199
transform 1 0 228 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1711653199
transform 1 0 164 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1711653199
transform 1 0 164 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1711653199
transform 1 0 132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1711653199
transform 1 0 964 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_1551
timestamp 1711653199
transform 1 0 940 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1552
timestamp 1711653199
transform 1 0 892 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1711653199
transform 1 0 868 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1711653199
transform 1 0 1036 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1711653199
transform 1 0 1020 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1711653199
transform 1 0 1556 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1711653199
transform 1 0 1556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1711653199
transform 1 0 932 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1711653199
transform 1 0 932 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1711653199
transform 1 0 908 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1711653199
transform 1 0 908 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1711653199
transform 1 0 908 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1711653199
transform 1 0 908 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1711653199
transform 1 0 1124 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1711653199
transform 1 0 1060 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1711653199
transform 1 0 1052 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1711653199
transform 1 0 1036 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1711653199
transform 1 0 1116 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1711653199
transform 1 0 1068 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1711653199
transform 1 0 1060 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1711653199
transform 1 0 1868 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1572
timestamp 1711653199
transform 1 0 1804 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1711653199
transform 1 0 1756 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1574
timestamp 1711653199
transform 1 0 1692 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1711653199
transform 1 0 1548 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1711653199
transform 1 0 1524 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1711653199
transform 1 0 1428 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1711653199
transform 1 0 1140 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1711653199
transform 1 0 1108 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1711653199
transform 1 0 1084 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1711653199
transform 1 0 1900 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1711653199
transform 1 0 1860 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1711653199
transform 1 0 1796 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1584
timestamp 1711653199
transform 1 0 1580 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1711653199
transform 1 0 1540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1711653199
transform 1 0 2284 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1711653199
transform 1 0 2252 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1711653199
transform 1 0 2236 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1589
timestamp 1711653199
transform 1 0 2236 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1711653199
transform 1 0 2124 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1711653199
transform 1 0 2068 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1592
timestamp 1711653199
transform 1 0 1196 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1711653199
transform 1 0 1196 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1711653199
transform 1 0 1188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1711653199
transform 1 0 1316 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_1596
timestamp 1711653199
transform 1 0 1316 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1711653199
transform 1 0 1196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1598
timestamp 1711653199
transform 1 0 1196 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_1599
timestamp 1711653199
transform 1 0 2420 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1711653199
transform 1 0 2276 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1711653199
transform 1 0 2156 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1711653199
transform 1 0 2108 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_1603
timestamp 1711653199
transform 1 0 1988 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1604
timestamp 1711653199
transform 1 0 1660 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1711653199
transform 1 0 1436 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1711653199
transform 1 0 3028 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1711653199
transform 1 0 2972 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1711653199
transform 1 0 2940 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1711653199
transform 1 0 3036 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1711653199
transform 1 0 3036 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_1611
timestamp 1711653199
transform 1 0 3332 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1711653199
transform 1 0 3316 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1711653199
transform 1 0 3364 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1711653199
transform 1 0 3364 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1711653199
transform 1 0 3308 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1616
timestamp 1711653199
transform 1 0 3284 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1617
timestamp 1711653199
transform 1 0 3252 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1711653199
transform 1 0 3372 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1711653199
transform 1 0 3308 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_1620
timestamp 1711653199
transform 1 0 3292 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1711653199
transform 1 0 3380 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1622
timestamp 1711653199
transform 1 0 3356 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1623
timestamp 1711653199
transform 1 0 3268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1711653199
transform 1 0 3356 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1711653199
transform 1 0 3356 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1711653199
transform 1 0 3332 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1711653199
transform 1 0 3380 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1711653199
transform 1 0 3324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1711653199
transform 1 0 3300 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1711653199
transform 1 0 3036 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1631
timestamp 1711653199
transform 1 0 3036 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1632
timestamp 1711653199
transform 1 0 2948 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1711653199
transform 1 0 2868 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1711653199
transform 1 0 2500 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1711653199
transform 1 0 2492 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1711653199
transform 1 0 2396 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1711653199
transform 1 0 2372 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1711653199
transform 1 0 2372 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1639
timestamp 1711653199
transform 1 0 2324 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1711653199
transform 1 0 2620 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1711653199
transform 1 0 2620 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1711653199
transform 1 0 2556 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1711653199
transform 1 0 2444 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1711653199
transform 1 0 2364 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1711653199
transform 1 0 2284 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1711653199
transform 1 0 2284 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1647
timestamp 1711653199
transform 1 0 2220 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1648
timestamp 1711653199
transform 1 0 2780 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1649
timestamp 1711653199
transform 1 0 2756 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1711653199
transform 1 0 2724 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1651
timestamp 1711653199
transform 1 0 2772 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1711653199
transform 1 0 2740 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1711653199
transform 1 0 2724 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1711653199
transform 1 0 2812 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1711653199
transform 1 0 2804 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1711653199
transform 1 0 2972 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1711653199
transform 1 0 2828 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1658
timestamp 1711653199
transform 1 0 2828 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1711653199
transform 1 0 1892 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1711653199
transform 1 0 1764 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1711653199
transform 1 0 1660 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1711653199
transform 1 0 1532 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1663
timestamp 1711653199
transform 1 0 1396 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1711653199
transform 1 0 1292 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1711653199
transform 1 0 1156 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1711653199
transform 1 0 1020 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1667
timestamp 1711653199
transform 1 0 876 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1711653199
transform 1 0 580 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1669
timestamp 1711653199
transform 1 0 468 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1670
timestamp 1711653199
transform 1 0 316 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1671
timestamp 1711653199
transform 1 0 316 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1672
timestamp 1711653199
transform 1 0 3204 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1673
timestamp 1711653199
transform 1 0 2820 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1711653199
transform 1 0 2732 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1711653199
transform 1 0 2612 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1711653199
transform 1 0 1884 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1711653199
transform 1 0 1716 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1711653199
transform 1 0 1500 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1679
timestamp 1711653199
transform 1 0 1268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1711653199
transform 1 0 788 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1711653199
transform 1 0 564 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1711653199
transform 1 0 420 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1711653199
transform 1 0 308 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1711653199
transform 1 0 276 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1711653199
transform 1 0 172 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1711653199
transform 1 0 172 0 1 3085
box -2 -2 2 2
use M2_M1  M2_M1_1687
timestamp 1711653199
transform 1 0 92 0 1 3085
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1711653199
transform 1 0 92 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1711653199
transform 1 0 92 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1711653199
transform 1 0 3316 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1711653199
transform 1 0 3316 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1692
timestamp 1711653199
transform 1 0 3268 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1711653199
transform 1 0 3220 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1711653199
transform 1 0 3004 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1711653199
transform 1 0 3004 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1711653199
transform 1 0 2980 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1711653199
transform 1 0 2812 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1711653199
transform 1 0 2748 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1711653199
transform 1 0 2644 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1700
timestamp 1711653199
transform 1 0 2596 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1701
timestamp 1711653199
transform 1 0 2564 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1711653199
transform 1 0 2500 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1711653199
transform 1 0 2468 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1704
timestamp 1711653199
transform 1 0 2452 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1705
timestamp 1711653199
transform 1 0 2444 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1711653199
transform 1 0 3316 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1711653199
transform 1 0 3308 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1711653199
transform 1 0 3092 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1711653199
transform 1 0 2900 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1710
timestamp 1711653199
transform 1 0 2900 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1711653199
transform 1 0 2804 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1712
timestamp 1711653199
transform 1 0 2716 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1711653199
transform 1 0 2508 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1711653199
transform 1 0 2372 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1711653199
transform 1 0 2276 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1711653199
transform 1 0 2172 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1711653199
transform 1 0 2076 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1711653199
transform 1 0 1972 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1711653199
transform 1 0 1900 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1720
timestamp 1711653199
transform 1 0 1924 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1711653199
transform 1 0 1852 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1711653199
transform 1 0 1812 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1711653199
transform 1 0 1708 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1711653199
transform 1 0 1572 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1725
timestamp 1711653199
transform 1 0 1468 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1711653199
transform 1 0 1300 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1711653199
transform 1 0 1004 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1711653199
transform 1 0 820 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1711653199
transform 1 0 692 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1711653199
transform 1 0 580 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1711653199
transform 1 0 428 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1711653199
transform 1 0 380 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1711653199
transform 1 0 276 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1711653199
transform 1 0 1964 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1711653199
transform 1 0 1860 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1711653199
transform 1 0 1828 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1711653199
transform 1 0 1780 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1711653199
transform 1 0 1724 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1711653199
transform 1 0 1508 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1711653199
transform 1 0 980 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1711653199
transform 1 0 732 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1742
timestamp 1711653199
transform 1 0 420 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1711653199
transform 1 0 340 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1711653199
transform 1 0 204 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1711653199
transform 1 0 92 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1711653199
transform 1 0 92 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1711653199
transform 1 0 92 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1748
timestamp 1711653199
transform 1 0 2556 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1711653199
transform 1 0 2556 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1711653199
transform 1 0 2444 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1711653199
transform 1 0 2340 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1711653199
transform 1 0 2300 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1753
timestamp 1711653199
transform 1 0 2236 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1711653199
transform 1 0 2196 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1711653199
transform 1 0 2188 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1711653199
transform 1 0 2036 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1711653199
transform 1 0 1628 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1711653199
transform 1 0 1516 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1711653199
transform 1 0 1476 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1711653199
transform 1 0 1412 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1711653199
transform 1 0 1364 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1711653199
transform 1 0 1244 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1711653199
transform 1 0 1156 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1711653199
transform 1 0 1044 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1711653199
transform 1 0 844 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1711653199
transform 1 0 812 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1767
timestamp 1711653199
transform 1 0 692 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1711653199
transform 1 0 580 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1711653199
transform 1 0 524 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1711653199
transform 1 0 460 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1711653199
transform 1 0 412 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1711653199
transform 1 0 308 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1711653199
transform 1 0 196 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1711653199
transform 1 0 92 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1711653199
transform 1 0 92 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1711653199
transform 1 0 3196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1711653199
transform 1 0 3164 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1711653199
transform 1 0 3068 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1711653199
transform 1 0 2980 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1711653199
transform 1 0 2876 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_1781
timestamp 1711653199
transform 1 0 2868 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1711653199
transform 1 0 2844 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1711653199
transform 1 0 2140 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1711653199
transform 1 0 2036 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1711653199
transform 1 0 1932 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1711653199
transform 1 0 1788 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1711653199
transform 1 0 1516 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1711653199
transform 1 0 1476 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1711653199
transform 1 0 1356 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1711653199
transform 1 0 1860 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1711653199
transform 1 0 1812 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1711653199
transform 1 0 1812 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1793
timestamp 1711653199
transform 1 0 1804 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1711653199
transform 1 0 1780 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1711653199
transform 1 0 1460 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1711653199
transform 1 0 1452 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1711653199
transform 1 0 1228 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1711653199
transform 1 0 2612 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1711653199
transform 1 0 2588 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1711653199
transform 1 0 2572 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1711653199
transform 1 0 2484 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1711653199
transform 1 0 3292 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1711653199
transform 1 0 3060 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1711653199
transform 1 0 2932 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1711653199
transform 1 0 2924 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1711653199
transform 1 0 2628 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1711653199
transform 1 0 2596 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1711653199
transform 1 0 2764 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1711653199
transform 1 0 2660 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1711653199
transform 1 0 2604 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1711653199
transform 1 0 2604 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1711653199
transform 1 0 2524 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1711653199
transform 1 0 2460 0 1 2785
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1711653199
transform 1 0 3268 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1711653199
transform 1 0 3052 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1711653199
transform 1 0 3012 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1711653199
transform 1 0 2988 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1711653199
transform 1 0 2940 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1711653199
transform 1 0 2860 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1711653199
transform 1 0 2740 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1711653199
transform 1 0 2564 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1822
timestamp 1711653199
transform 1 0 2028 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1711653199
transform 1 0 2012 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_1824
timestamp 1711653199
transform 1 0 1796 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1711653199
transform 1 0 1780 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1711653199
transform 1 0 1484 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1711653199
transform 1 0 932 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1711653199
transform 1 0 668 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1711653199
transform 1 0 516 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1830
timestamp 1711653199
transform 1 0 364 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1711653199
transform 1 0 348 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1711653199
transform 1 0 260 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1711653199
transform 1 0 228 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1834
timestamp 1711653199
transform 1 0 228 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1711653199
transform 1 0 212 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1711653199
transform 1 0 204 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1711653199
transform 1 0 196 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1711653199
transform 1 0 2124 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1711653199
transform 1 0 2060 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1711653199
transform 1 0 2036 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1711653199
transform 1 0 1908 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1842
timestamp 1711653199
transform 1 0 1836 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1711653199
transform 1 0 1740 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1844
timestamp 1711653199
transform 1 0 1948 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1845
timestamp 1711653199
transform 1 0 1852 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1711653199
transform 1 0 1668 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1711653199
transform 1 0 1636 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1711653199
transform 1 0 1756 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1711653199
transform 1 0 1388 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1850
timestamp 1711653199
transform 1 0 1324 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1851
timestamp 1711653199
transform 1 0 932 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1852
timestamp 1711653199
transform 1 0 828 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1853
timestamp 1711653199
transform 1 0 764 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1711653199
transform 1 0 572 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1711653199
transform 1 0 548 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1711653199
transform 1 0 2348 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1711653199
transform 1 0 1940 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1858
timestamp 1711653199
transform 1 0 476 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1711653199
transform 1 0 436 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1711653199
transform 1 0 404 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1711653199
transform 1 0 292 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1711653199
transform 1 0 252 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1863
timestamp 1711653199
transform 1 0 212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1711653199
transform 1 0 124 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1711653199
transform 1 0 2148 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1711653199
transform 1 0 2052 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1867
timestamp 1711653199
transform 1 0 1868 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1868
timestamp 1711653199
transform 1 0 1612 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1869
timestamp 1711653199
transform 1 0 1260 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1711653199
transform 1 0 1156 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1871
timestamp 1711653199
transform 1 0 1132 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1711653199
transform 1 0 1092 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1711653199
transform 1 0 2108 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1711653199
transform 1 0 2084 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1711653199
transform 1 0 2084 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1711653199
transform 1 0 2652 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1711653199
transform 1 0 2532 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1878
timestamp 1711653199
transform 1 0 2284 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1879
timestamp 1711653199
transform 1 0 2156 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1880
timestamp 1711653199
transform 1 0 1892 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1711653199
transform 1 0 1860 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1882
timestamp 1711653199
transform 1 0 1684 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1711653199
transform 1 0 1588 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1884
timestamp 1711653199
transform 1 0 2180 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_1885
timestamp 1711653199
transform 1 0 2180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1711653199
transform 1 0 2140 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1711653199
transform 1 0 2140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1888
timestamp 1711653199
transform 1 0 2100 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1889
timestamp 1711653199
transform 1 0 1988 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1890
timestamp 1711653199
transform 1 0 1908 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1711653199
transform 1 0 1652 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1711653199
transform 1 0 1636 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1893
timestamp 1711653199
transform 1 0 1428 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1894
timestamp 1711653199
transform 1 0 1364 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1895
timestamp 1711653199
transform 1 0 1300 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1896
timestamp 1711653199
transform 1 0 1212 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1711653199
transform 1 0 1148 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1711653199
transform 1 0 1124 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1711653199
transform 1 0 948 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1900
timestamp 1711653199
transform 1 0 884 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1711653199
transform 1 0 820 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1902
timestamp 1711653199
transform 1 0 628 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1903
timestamp 1711653199
transform 1 0 372 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_1904
timestamp 1711653199
transform 1 0 268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1905
timestamp 1711653199
transform 1 0 244 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1711653199
transform 1 0 2684 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1711653199
transform 1 0 2668 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1908
timestamp 1711653199
transform 1 0 2604 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1711653199
transform 1 0 2364 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1711653199
transform 1 0 2724 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1911
timestamp 1711653199
transform 1 0 2476 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_1912
timestamp 1711653199
transform 1 0 2236 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1711653199
transform 1 0 1980 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1914
timestamp 1711653199
transform 1 0 2348 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1915
timestamp 1711653199
transform 1 0 2332 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1916
timestamp 1711653199
transform 1 0 2308 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_1917
timestamp 1711653199
transform 1 0 2172 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1918
timestamp 1711653199
transform 1 0 2092 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1919
timestamp 1711653199
transform 1 0 1812 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1920
timestamp 1711653199
transform 1 0 1724 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1921
timestamp 1711653199
transform 1 0 1684 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1711653199
transform 1 0 1676 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1711653199
transform 1 0 1652 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_1924
timestamp 1711653199
transform 1 0 1564 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1711653199
transform 1 0 1556 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1926
timestamp 1711653199
transform 1 0 1460 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1711653199
transform 1 0 1372 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1711653199
transform 1 0 1220 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1711653199
transform 1 0 1100 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1711653199
transform 1 0 1020 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1711653199
transform 1 0 940 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1932
timestamp 1711653199
transform 1 0 724 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1711653199
transform 1 0 628 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1711653199
transform 1 0 604 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1711653199
transform 1 0 596 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1711653199
transform 1 0 564 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1711653199
transform 1 0 556 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1711653199
transform 1 0 524 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1711653199
transform 1 0 508 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1711653199
transform 1 0 492 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1711653199
transform 1 0 468 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1711653199
transform 1 0 444 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1711653199
transform 1 0 428 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1711653199
transform 1 0 2316 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1711653199
transform 1 0 2204 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1711653199
transform 1 0 2148 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1711653199
transform 1 0 2036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1711653199
transform 1 0 1956 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1711653199
transform 1 0 1836 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1711653199
transform 1 0 1820 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1711653199
transform 1 0 1708 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1711653199
transform 1 0 1700 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1711653199
transform 1 0 1588 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1711653199
transform 1 0 1564 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1711653199
transform 1 0 1436 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1711653199
transform 1 0 1388 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1711653199
transform 1 0 1308 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1711653199
transform 1 0 1140 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1711653199
transform 1 0 1020 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1711653199
transform 1 0 916 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1711653199
transform 1 0 908 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1962
timestamp 1711653199
transform 1 0 692 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1711653199
transform 1 0 676 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1711653199
transform 1 0 532 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1711653199
transform 1 0 492 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1711653199
transform 1 0 412 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1711653199
transform 1 0 364 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_1968
timestamp 1711653199
transform 1 0 332 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1711653199
transform 1 0 228 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1711653199
transform 1 0 220 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1711653199
transform 1 0 220 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1711653199
transform 1 0 204 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_1973
timestamp 1711653199
transform 1 0 3188 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1711653199
transform 1 0 3156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_1975
timestamp 1711653199
transform 1 0 3068 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1711653199
transform 1 0 3060 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1711653199
transform 1 0 2684 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1711653199
transform 1 0 2252 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1711653199
transform 1 0 3012 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1980
timestamp 1711653199
transform 1 0 2996 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1711653199
transform 1 0 2916 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1711653199
transform 1 0 2884 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1711653199
transform 1 0 2868 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1711653199
transform 1 0 3300 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1711653199
transform 1 0 3300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1711653199
transform 1 0 3100 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1711653199
transform 1 0 2644 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1711653199
transform 1 0 2308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1711653199
transform 1 0 2260 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1711653199
transform 1 0 2244 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_1991
timestamp 1711653199
transform 1 0 2180 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1711653199
transform 1 0 2124 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1711653199
transform 1 0 2124 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1711653199
transform 1 0 2100 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1711653199
transform 1 0 2068 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1711653199
transform 1 0 2028 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1711653199
transform 1 0 2028 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1711653199
transform 1 0 1948 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1711653199
transform 1 0 1628 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1711653199
transform 1 0 1580 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1711653199
transform 1 0 1388 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1711653199
transform 1 0 1220 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1711653199
transform 1 0 1132 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1711653199
transform 1 0 1116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1711653199
transform 1 0 1100 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1711653199
transform 1 0 1100 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1711653199
transform 1 0 980 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1711653199
transform 1 0 876 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1711653199
transform 1 0 844 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1711653199
transform 1 0 700 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1711653199
transform 1 0 684 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1711653199
transform 1 0 684 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1711653199
transform 1 0 668 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1711653199
transform 1 0 612 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1711653199
transform 1 0 612 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1711653199
transform 1 0 388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1711653199
transform 1 0 244 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1711653199
transform 1 0 236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1711653199
transform 1 0 220 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1711653199
transform 1 0 180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1711653199
transform 1 0 172 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2022
timestamp 1711653199
transform 1 0 3028 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1711653199
transform 1 0 2988 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1711653199
transform 1 0 2916 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1711653199
transform 1 0 2748 0 1 1785
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1711653199
transform 1 0 2580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1711653199
transform 1 0 2548 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1711653199
transform 1 0 2444 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1711653199
transform 1 0 2276 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1711653199
transform 1 0 2236 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1711653199
transform 1 0 2140 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1711653199
transform 1 0 3300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2033
timestamp 1711653199
transform 1 0 3300 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1711653199
transform 1 0 3260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1711653199
transform 1 0 3164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1711653199
transform 1 0 2940 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1711653199
transform 1 0 2708 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1711653199
transform 1 0 2564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1711653199
transform 1 0 2012 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1711653199
transform 1 0 1964 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1711653199
transform 1 0 1932 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1711653199
transform 1 0 1908 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1711653199
transform 1 0 1732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1711653199
transform 1 0 1692 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1711653199
transform 1 0 1652 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1711653199
transform 1 0 1524 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1711653199
transform 1 0 1500 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1711653199
transform 1 0 1428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1711653199
transform 1 0 1284 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1711653199
transform 1 0 1036 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1711653199
transform 1 0 988 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1711653199
transform 1 0 796 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1711653199
transform 1 0 748 0 1 1445
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1711653199
transform 1 0 652 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1711653199
transform 1 0 652 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1711653199
transform 1 0 532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1711653199
transform 1 0 380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1711653199
transform 1 0 372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1711653199
transform 1 0 324 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1711653199
transform 1 0 244 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1711653199
transform 1 0 196 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1711653199
transform 1 0 3188 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2063
timestamp 1711653199
transform 1 0 3164 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1711653199
transform 1 0 2804 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_2065
timestamp 1711653199
transform 1 0 3188 0 1 2055
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1711653199
transform 1 0 3188 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1711653199
transform 1 0 3164 0 1 2055
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1711653199
transform 1 0 3140 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1711653199
transform 1 0 2884 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1711653199
transform 1 0 2700 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1711653199
transform 1 0 2684 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2072
timestamp 1711653199
transform 1 0 3180 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2073
timestamp 1711653199
transform 1 0 3180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1711653199
transform 1 0 3132 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1711653199
transform 1 0 2636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1711653199
transform 1 0 2516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1711653199
transform 1 0 1700 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1711653199
transform 1 0 1628 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_2079
timestamp 1711653199
transform 1 0 1348 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1711653199
transform 1 0 1228 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1711653199
transform 1 0 996 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1711653199
transform 1 0 908 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2083
timestamp 1711653199
transform 1 0 764 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1711653199
transform 1 0 684 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1711653199
transform 1 0 484 0 1 1455
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1711653199
transform 1 0 348 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1711653199
transform 1 0 292 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1711653199
transform 1 0 3260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1711653199
transform 1 0 3236 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1711653199
transform 1 0 3028 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1711653199
transform 1 0 2956 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1711653199
transform 1 0 2372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1711653199
transform 1 0 2284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1711653199
transform 1 0 2116 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1711653199
transform 1 0 1900 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1711653199
transform 1 0 1868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1711653199
transform 1 0 1844 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1711653199
transform 1 0 1788 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2099
timestamp 1711653199
transform 1 0 1572 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2100
timestamp 1711653199
transform 1 0 620 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1711653199
transform 1 0 604 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1711653199
transform 1 0 604 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1711653199
transform 1 0 332 0 1 1445
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1711653199
transform 1 0 204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1711653199
transform 1 0 156 0 1 1695
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1711653199
transform 1 0 3140 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1711653199
transform 1 0 3108 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2108
timestamp 1711653199
transform 1 0 3116 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2109
timestamp 1711653199
transform 1 0 2492 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2110
timestamp 1711653199
transform 1 0 2396 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1711653199
transform 1 0 2380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1711653199
transform 1 0 3260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1711653199
transform 1 0 3220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2114
timestamp 1711653199
transform 1 0 3108 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1711653199
transform 1 0 3044 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1711653199
transform 1 0 2972 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2117
timestamp 1711653199
transform 1 0 2956 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1711653199
transform 1 0 2748 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2119
timestamp 1711653199
transform 1 0 2508 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1711653199
transform 1 0 2460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1711653199
transform 1 0 2292 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1711653199
transform 1 0 2204 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2123
timestamp 1711653199
transform 1 0 1996 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1711653199
transform 1 0 1996 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1711653199
transform 1 0 1924 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1711653199
transform 1 0 1788 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1711653199
transform 1 0 1348 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1711653199
transform 1 0 1316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2129
timestamp 1711653199
transform 1 0 1116 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1711653199
transform 1 0 1100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1711653199
transform 1 0 780 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1711653199
transform 1 0 588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1711653199
transform 1 0 484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1711653199
transform 1 0 436 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1711653199
transform 1 0 332 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1711653199
transform 1 0 180 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2137
timestamp 1711653199
transform 1 0 172 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1711653199
transform 1 0 148 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2139
timestamp 1711653199
transform 1 0 140 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1711653199
transform 1 0 140 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1711653199
transform 1 0 2628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1711653199
transform 1 0 2612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1711653199
transform 1 0 2380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1711653199
transform 1 0 2252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2145
timestamp 1711653199
transform 1 0 2100 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2146
timestamp 1711653199
transform 1 0 1940 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2147
timestamp 1711653199
transform 1 0 1876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1711653199
transform 1 0 1724 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1711653199
transform 1 0 1252 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1711653199
transform 1 0 1052 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2151
timestamp 1711653199
transform 1 0 1020 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1711653199
transform 1 0 556 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1711653199
transform 1 0 420 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1711653199
transform 1 0 404 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1711653199
transform 1 0 3332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1711653199
transform 1 0 3316 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1711653199
transform 1 0 3124 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1711653199
transform 1 0 2796 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1711653199
transform 1 0 2348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2160
timestamp 1711653199
transform 1 0 1364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1711653199
transform 1 0 924 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1711653199
transform 1 0 636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1711653199
transform 1 0 412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1711653199
transform 1 0 372 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1711653199
transform 1 0 260 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1711653199
transform 1 0 252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1711653199
transform 1 0 172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1711653199
transform 1 0 140 0 1 695
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1711653199
transform 1 0 2972 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1711653199
transform 1 0 2876 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2171
timestamp 1711653199
transform 1 0 2836 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1711653199
transform 1 0 3156 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1711653199
transform 1 0 3116 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2174
timestamp 1711653199
transform 1 0 2948 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1711653199
transform 1 0 2860 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1711653199
transform 1 0 3300 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1711653199
transform 1 0 3204 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1711653199
transform 1 0 3132 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1711653199
transform 1 0 3100 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1711653199
transform 1 0 3068 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1711653199
transform 1 0 2924 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1711653199
transform 1 0 2916 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1711653199
transform 1 0 2732 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1711653199
transform 1 0 2732 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1711653199
transform 1 0 2476 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1711653199
transform 1 0 2428 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1711653199
transform 1 0 2284 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1711653199
transform 1 0 2252 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2189
timestamp 1711653199
transform 1 0 2188 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2190
timestamp 1711653199
transform 1 0 2188 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1711653199
transform 1 0 2172 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1711653199
transform 1 0 2052 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2193
timestamp 1711653199
transform 1 0 2028 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1711653199
transform 1 0 1804 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1711653199
transform 1 0 1764 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1711653199
transform 1 0 1676 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1711653199
transform 1 0 1580 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1711653199
transform 1 0 1564 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1711653199
transform 1 0 1420 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1711653199
transform 1 0 1348 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1711653199
transform 1 0 1172 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1711653199
transform 1 0 1124 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1711653199
transform 1 0 916 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1711653199
transform 1 0 540 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1711653199
transform 1 0 516 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2206
timestamp 1711653199
transform 1 0 516 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1711653199
transform 1 0 484 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1711653199
transform 1 0 444 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1711653199
transform 1 0 164 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1711653199
transform 1 0 124 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1711653199
transform 1 0 116 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2212
timestamp 1711653199
transform 1 0 108 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1711653199
transform 1 0 2996 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1711653199
transform 1 0 2892 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2215
timestamp 1711653199
transform 1 0 2884 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1711653199
transform 1 0 2852 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1711653199
transform 1 0 2244 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1711653199
transform 1 0 1916 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1711653199
transform 1 0 1852 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1711653199
transform 1 0 1772 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2221
timestamp 1711653199
transform 1 0 1724 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1711653199
transform 1 0 1556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1711653199
transform 1 0 1396 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1711653199
transform 1 0 1220 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1711653199
transform 1 0 1084 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1711653199
transform 1 0 948 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1711653199
transform 1 0 828 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1711653199
transform 1 0 3356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2229
timestamp 1711653199
transform 1 0 3260 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2230
timestamp 1711653199
transform 1 0 3132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2231
timestamp 1711653199
transform 1 0 3100 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_2232
timestamp 1711653199
transform 1 0 2860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2233
timestamp 1711653199
transform 1 0 2220 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1711653199
transform 1 0 2212 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1711653199
transform 1 0 2196 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1711653199
transform 1 0 1820 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1711653199
transform 1 0 1748 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2238
timestamp 1711653199
transform 1 0 1700 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1711653199
transform 1 0 1500 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2240
timestamp 1711653199
transform 1 0 1356 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1711653199
transform 1 0 1180 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1711653199
transform 1 0 1100 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2243
timestamp 1711653199
transform 1 0 788 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2244
timestamp 1711653199
transform 1 0 404 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1711653199
transform 1 0 332 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1711653199
transform 1 0 180 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1711653199
transform 1 0 3092 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1711653199
transform 1 0 2980 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1711653199
transform 1 0 2956 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1711653199
transform 1 0 2204 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1711653199
transform 1 0 2036 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1711653199
transform 1 0 1988 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1711653199
transform 1 0 1876 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2254
timestamp 1711653199
transform 1 0 1660 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1711653199
transform 1 0 1452 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1711653199
transform 1 0 1260 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1711653199
transform 1 0 1100 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1711653199
transform 1 0 460 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1711653199
transform 1 0 420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1711653199
transform 1 0 340 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1711653199
transform 1 0 236 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1711653199
transform 1 0 188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1711653199
transform 1 0 100 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1711653199
transform 1 0 2588 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1711653199
transform 1 0 2444 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1711653199
transform 1 0 2404 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1711653199
transform 1 0 2276 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1711653199
transform 1 0 2244 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1711653199
transform 1 0 1620 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1711653199
transform 1 0 1420 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1711653199
transform 1 0 1364 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1711653199
transform 1 0 1308 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1711653199
transform 1 0 956 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2274
timestamp 1711653199
transform 1 0 900 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1711653199
transform 1 0 620 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1711653199
transform 1 0 564 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1711653199
transform 1 0 532 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1711653199
transform 1 0 3148 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1711653199
transform 1 0 3132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1711653199
transform 1 0 3092 0 1 2485
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1711653199
transform 1 0 3076 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1711653199
transform 1 0 2940 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1711653199
transform 1 0 2812 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1711653199
transform 1 0 2772 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1711653199
transform 1 0 2652 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1711653199
transform 1 0 2436 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1711653199
transform 1 0 2404 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1711653199
transform 1 0 2404 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1711653199
transform 1 0 2364 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1711653199
transform 1 0 2308 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1711653199
transform 1 0 2156 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1711653199
transform 1 0 2820 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1711653199
transform 1 0 2820 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1711653199
transform 1 0 2804 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1711653199
transform 1 0 2180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1711653199
transform 1 0 2092 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2297
timestamp 1711653199
transform 1 0 1852 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1711653199
transform 1 0 1700 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2299
timestamp 1711653199
transform 1 0 1628 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2300
timestamp 1711653199
transform 1 0 1044 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1711653199
transform 1 0 1004 0 1 1095
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1711653199
transform 1 0 1004 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1711653199
transform 1 0 996 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1711653199
transform 1 0 964 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2305
timestamp 1711653199
transform 1 0 844 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1711653199
transform 1 0 796 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1711653199
transform 1 0 740 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2308
timestamp 1711653199
transform 1 0 652 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1711653199
transform 1 0 644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1711653199
transform 1 0 2852 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1711653199
transform 1 0 2852 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1711653199
transform 1 0 2828 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1711653199
transform 1 0 2596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1711653199
transform 1 0 2548 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1711653199
transform 1 0 2468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1711653199
transform 1 0 2380 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1711653199
transform 1 0 1884 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1711653199
transform 1 0 1836 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2319
timestamp 1711653199
transform 1 0 1796 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1711653199
transform 1 0 1196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2321
timestamp 1711653199
transform 1 0 1180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1711653199
transform 1 0 996 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1711653199
transform 1 0 996 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1711653199
transform 1 0 964 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1711653199
transform 1 0 964 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1711653199
transform 1 0 780 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1711653199
transform 1 0 764 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1711653199
transform 1 0 700 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1711653199
transform 1 0 676 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2330
timestamp 1711653199
transform 1 0 676 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1711653199
transform 1 0 3140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2332
timestamp 1711653199
transform 1 0 3108 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1711653199
transform 1 0 3100 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1711653199
transform 1 0 3052 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1711653199
transform 1 0 2252 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1711653199
transform 1 0 1972 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2337
timestamp 1711653199
transform 1 0 1804 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1711653199
transform 1 0 1724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2339
timestamp 1711653199
transform 1 0 1620 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_2340
timestamp 1711653199
transform 1 0 1340 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2341
timestamp 1711653199
transform 1 0 812 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1711653199
transform 1 0 804 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1711653199
transform 1 0 780 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1711653199
transform 1 0 668 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2345
timestamp 1711653199
transform 1 0 524 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1711653199
transform 1 0 436 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2347
timestamp 1711653199
transform 1 0 348 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1711653199
transform 1 0 348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1711653199
transform 1 0 2204 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1711653199
transform 1 0 2148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1711653199
transform 1 0 2148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2352
timestamp 1711653199
transform 1 0 1780 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1711653199
transform 1 0 1084 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1711653199
transform 1 0 1028 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1711653199
transform 1 0 972 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2356
timestamp 1711653199
transform 1 0 748 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2357
timestamp 1711653199
transform 1 0 676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1711653199
transform 1 0 620 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2359
timestamp 1711653199
transform 1 0 564 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2360
timestamp 1711653199
transform 1 0 3284 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1711653199
transform 1 0 3284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1711653199
transform 1 0 3060 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1711653199
transform 1 0 2772 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2364
timestamp 1711653199
transform 1 0 2412 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1711653199
transform 1 0 1748 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1711653199
transform 1 0 1604 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2367
timestamp 1711653199
transform 1 0 1540 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1711653199
transform 1 0 1484 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1711653199
transform 1 0 1308 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1711653199
transform 1 0 812 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1711653199
transform 1 0 556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1711653199
transform 1 0 284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1711653199
transform 1 0 212 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2374
timestamp 1711653199
transform 1 0 180 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1711653199
transform 1 0 100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1711653199
transform 1 0 68 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1711653199
transform 1 0 2524 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1711653199
transform 1 0 2508 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1711653199
transform 1 0 2508 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1711653199
transform 1 0 2468 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1711653199
transform 1 0 2332 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1711653199
transform 1 0 1708 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1711653199
transform 1 0 1596 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1711653199
transform 1 0 1356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2385
timestamp 1711653199
transform 1 0 1132 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2386
timestamp 1711653199
transform 1 0 1116 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1711653199
transform 1 0 1116 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1711653199
transform 1 0 780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1711653199
transform 1 0 740 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2390
timestamp 1711653199
transform 1 0 596 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2391
timestamp 1711653199
transform 1 0 588 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1711653199
transform 1 0 324 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1711653199
transform 1 0 308 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1711653199
transform 1 0 292 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1711653199
transform 1 0 1268 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2396
timestamp 1711653199
transform 1 0 1108 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1711653199
transform 1 0 1052 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1711653199
transform 1 0 956 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2399
timestamp 1711653199
transform 1 0 852 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1711653199
transform 1 0 852 0 1 1285
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1711653199
transform 1 0 852 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1711653199
transform 1 0 836 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1711653199
transform 1 0 836 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1711653199
transform 1 0 836 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1711653199
transform 1 0 828 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_2406
timestamp 1711653199
transform 1 0 820 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1711653199
transform 1 0 668 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_2408
timestamp 1711653199
transform 1 0 660 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1711653199
transform 1 0 660 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1711653199
transform 1 0 660 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1711653199
transform 1 0 452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1711653199
transform 1 0 268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2413
timestamp 1711653199
transform 1 0 260 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1711653199
transform 1 0 3092 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1711653199
transform 1 0 3036 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1711653199
transform 1 0 2972 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2417
timestamp 1711653199
transform 1 0 3308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1711653199
transform 1 0 3196 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_2419
timestamp 1711653199
transform 1 0 3172 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1711653199
transform 1 0 3172 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1711653199
transform 1 0 3252 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1711653199
transform 1 0 2956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2423
timestamp 1711653199
transform 1 0 2396 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1711653199
transform 1 0 3004 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2425
timestamp 1711653199
transform 1 0 2908 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1711653199
transform 1 0 2732 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1711653199
transform 1 0 2196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1711653199
transform 1 0 2172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1711653199
transform 1 0 2036 0 1 2155
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1711653199
transform 1 0 1244 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_2431
timestamp 1711653199
transform 1 0 1204 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_2432
timestamp 1711653199
transform 1 0 1148 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1711653199
transform 1 0 996 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1711653199
transform 1 0 2868 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1711653199
transform 1 0 2844 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1711653199
transform 1 0 2780 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1711653199
transform 1 0 2644 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1711653199
transform 1 0 2564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1711653199
transform 1 0 2244 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1711653199
transform 1 0 1996 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1711653199
transform 1 0 1812 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1711653199
transform 1 0 1812 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1711653199
transform 1 0 2756 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1711653199
transform 1 0 2692 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1711653199
transform 1 0 2668 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1711653199
transform 1 0 3156 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1711653199
transform 1 0 3100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1711653199
transform 1 0 3084 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1711653199
transform 1 0 3084 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1711653199
transform 1 0 3068 0 1 1045
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1711653199
transform 1 0 3068 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1711653199
transform 1 0 3068 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1711653199
transform 1 0 3012 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2454
timestamp 1711653199
transform 1 0 2956 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1711653199
transform 1 0 2932 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1711653199
transform 1 0 2956 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1711653199
transform 1 0 2812 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1711653199
transform 1 0 2748 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1711653199
transform 1 0 2268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1711653199
transform 1 0 2900 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1711653199
transform 1 0 2788 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1711653199
transform 1 0 2788 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1711653199
transform 1 0 2084 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2464
timestamp 1711653199
transform 1 0 2036 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1711653199
transform 1 0 2012 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1711653199
transform 1 0 1284 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1711653199
transform 1 0 1244 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1711653199
transform 1 0 892 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2469
timestamp 1711653199
transform 1 0 828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1711653199
transform 1 0 764 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1711653199
transform 1 0 716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1711653199
transform 1 0 2620 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1711653199
transform 1 0 2308 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1711653199
transform 1 0 2836 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1711653199
transform 1 0 2748 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2476
timestamp 1711653199
transform 1 0 2700 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2477
timestamp 1711653199
transform 1 0 2732 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1711653199
transform 1 0 2700 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1711653199
transform 1 0 3396 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1711653199
transform 1 0 3356 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1711653199
transform 1 0 3348 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_2482
timestamp 1711653199
transform 1 0 3316 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2483
timestamp 1711653199
transform 1 0 2820 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2484
timestamp 1711653199
transform 1 0 2788 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1711653199
transform 1 0 2764 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1711653199
transform 1 0 324 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1711653199
transform 1 0 292 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1711653199
transform 1 0 260 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1711653199
transform 1 0 148 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1711653199
transform 1 0 92 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1711653199
transform 1 0 2812 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1711653199
transform 1 0 2724 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1711653199
transform 1 0 2636 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2494
timestamp 1711653199
transform 1 0 2636 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1711653199
transform 1 0 2188 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1711653199
transform 1 0 2156 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1711653199
transform 1 0 2028 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1711653199
transform 1 0 1748 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2499
timestamp 1711653199
transform 1 0 1132 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1711653199
transform 1 0 988 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1711653199
transform 1 0 988 0 1 1485
box -2 -2 2 2
use M2_M1  M2_M1_2502
timestamp 1711653199
transform 1 0 948 0 1 1485
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1711653199
transform 1 0 924 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2504
timestamp 1711653199
transform 1 0 3364 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1711653199
transform 1 0 3348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1711653199
transform 1 0 3300 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1711653199
transform 1 0 3292 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1711653199
transform 1 0 2964 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1711653199
transform 1 0 2884 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1711653199
transform 1 0 2820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1711653199
transform 1 0 2748 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1711653199
transform 1 0 3116 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1711653199
transform 1 0 3012 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1711653199
transform 1 0 2916 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1711653199
transform 1 0 2900 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1711653199
transform 1 0 2780 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1711653199
transform 1 0 2780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2518
timestamp 1711653199
transform 1 0 2772 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1711653199
transform 1 0 2708 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1711653199
transform 1 0 3164 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1711653199
transform 1 0 3052 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1711653199
transform 1 0 3132 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2523
timestamp 1711653199
transform 1 0 3052 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1711653199
transform 1 0 2932 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1711653199
transform 1 0 2860 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1711653199
transform 1 0 2764 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2527
timestamp 1711653199
transform 1 0 2692 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1711653199
transform 1 0 2732 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1711653199
transform 1 0 2644 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2530
timestamp 1711653199
transform 1 0 3340 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2531
timestamp 1711653199
transform 1 0 3340 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1711653199
transform 1 0 3324 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2533
timestamp 1711653199
transform 1 0 3268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1711653199
transform 1 0 3084 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1711653199
transform 1 0 3068 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1711653199
transform 1 0 3004 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1711653199
transform 1 0 2980 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1711653199
transform 1 0 2932 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1711653199
transform 1 0 2932 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1711653199
transform 1 0 2812 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1711653199
transform 1 0 3132 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1711653199
transform 1 0 3116 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2543
timestamp 1711653199
transform 1 0 3188 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1711653199
transform 1 0 3188 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1711653199
transform 1 0 2964 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2546
timestamp 1711653199
transform 1 0 2892 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1711653199
transform 1 0 2868 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1711653199
transform 1 0 2812 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1711653199
transform 1 0 2908 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1711653199
transform 1 0 2828 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1711653199
transform 1 0 3228 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1711653199
transform 1 0 3148 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2553
timestamp 1711653199
transform 1 0 3108 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1711653199
transform 1 0 3028 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_2555
timestamp 1711653199
transform 1 0 2436 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1711653199
transform 1 0 2284 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1711653199
transform 1 0 2468 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1711653199
transform 1 0 2388 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2559
timestamp 1711653199
transform 1 0 2388 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2560
timestamp 1711653199
transform 1 0 2348 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1711653199
transform 1 0 2356 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2562
timestamp 1711653199
transform 1 0 2236 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2563
timestamp 1711653199
transform 1 0 2468 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1711653199
transform 1 0 2436 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1711653199
transform 1 0 2676 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2566
timestamp 1711653199
transform 1 0 2604 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2567
timestamp 1711653199
transform 1 0 2612 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1711653199
transform 1 0 2596 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1711653199
transform 1 0 2300 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1711653199
transform 1 0 2076 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1711653199
transform 1 0 2276 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1711653199
transform 1 0 2244 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1711653199
transform 1 0 1540 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1711653199
transform 1 0 1420 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1711653199
transform 1 0 1660 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1711653199
transform 1 0 1652 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2577
timestamp 1711653199
transform 1 0 1388 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_2578
timestamp 1711653199
transform 1 0 1372 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1711653199
transform 1 0 1444 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2580
timestamp 1711653199
transform 1 0 1436 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1711653199
transform 1 0 716 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1711653199
transform 1 0 604 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1711653199
transform 1 0 652 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2584
timestamp 1711653199
transform 1 0 620 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1711653199
transform 1 0 948 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1711653199
transform 1 0 892 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2587
timestamp 1711653199
transform 1 0 980 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2588
timestamp 1711653199
transform 1 0 860 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2589
timestamp 1711653199
transform 1 0 556 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1711653199
transform 1 0 548 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1711653199
transform 1 0 452 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1711653199
transform 1 0 452 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1711653199
transform 1 0 508 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1711653199
transform 1 0 500 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2595
timestamp 1711653199
transform 1 0 132 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1711653199
transform 1 0 132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1711653199
transform 1 0 228 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1711653199
transform 1 0 124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1711653199
transform 1 0 260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2600
timestamp 1711653199
transform 1 0 244 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1711653199
transform 1 0 364 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1711653199
transform 1 0 356 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1711653199
transform 1 0 1140 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1711653199
transform 1 0 1092 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1711653199
transform 1 0 1316 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1711653199
transform 1 0 1204 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1711653199
transform 1 0 1476 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1711653199
transform 1 0 1404 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2609
timestamp 1711653199
transform 1 0 1684 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2610
timestamp 1711653199
transform 1 0 1564 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1711653199
transform 1 0 1932 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1711653199
transform 1 0 1836 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2613
timestamp 1711653199
transform 1 0 2028 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1711653199
transform 1 0 1980 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1711653199
transform 1 0 2092 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1711653199
transform 1 0 2084 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2617
timestamp 1711653199
transform 1 0 2180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_2618
timestamp 1711653199
transform 1 0 2180 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1711653199
transform 1 0 1748 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1711653199
transform 1 0 1724 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1711653199
transform 1 0 3228 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1711653199
transform 1 0 3204 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1711653199
transform 1 0 2996 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1711653199
transform 1 0 2876 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2625
timestamp 1711653199
transform 1 0 1828 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1711653199
transform 1 0 1644 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1711653199
transform 1 0 1564 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2628
timestamp 1711653199
transform 1 0 1556 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2629
timestamp 1711653199
transform 1 0 1356 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1711653199
transform 1 0 780 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2631
timestamp 1711653199
transform 1 0 636 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1711653199
transform 1 0 468 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2633
timestamp 1711653199
transform 1 0 276 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1711653199
transform 1 0 228 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2635
timestamp 1711653199
transform 1 0 220 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1711653199
transform 1 0 212 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1711653199
transform 1 0 3172 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2638
timestamp 1711653199
transform 1 0 3132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1711653199
transform 1 0 2964 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1711653199
transform 1 0 2732 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2641
timestamp 1711653199
transform 1 0 2284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1711653199
transform 1 0 2124 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1711653199
transform 1 0 1668 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1711653199
transform 1 0 1316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2645
timestamp 1711653199
transform 1 0 748 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2646
timestamp 1711653199
transform 1 0 700 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1711653199
transform 1 0 588 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1711653199
transform 1 0 388 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2649
timestamp 1711653199
transform 1 0 220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1711653199
transform 1 0 196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1711653199
transform 1 0 140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1711653199
transform 1 0 140 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1711653199
transform 1 0 1644 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1711653199
transform 1 0 1548 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1711653199
transform 1 0 1748 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1711653199
transform 1 0 1628 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1711653199
transform 1 0 3204 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1711653199
transform 1 0 3188 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1711653199
transform 1 0 3164 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1711653199
transform 1 0 3140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1711653199
transform 1 0 3100 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1711653199
transform 1 0 2908 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_2663
timestamp 1711653199
transform 1 0 2732 0 1 2385
box -2 -2 2 2
use M2_M1  M2_M1_2664
timestamp 1711653199
transform 1 0 2708 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1711653199
transform 1 0 3228 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_2666
timestamp 1711653199
transform 1 0 3140 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2667
timestamp 1711653199
transform 1 0 2452 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2668
timestamp 1711653199
transform 1 0 2388 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2669
timestamp 1711653199
transform 1 0 2356 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1711653199
transform 1 0 3332 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2671
timestamp 1711653199
transform 1 0 3284 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1711653199
transform 1 0 3356 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2673
timestamp 1711653199
transform 1 0 3340 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1711653199
transform 1 0 3244 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1711653199
transform 1 0 3220 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1711653199
transform 1 0 3164 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_2677
timestamp 1711653199
transform 1 0 3060 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1711653199
transform 1 0 3020 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2679
timestamp 1711653199
transform 1 0 2940 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1711653199
transform 1 0 2868 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1711653199
transform 1 0 2772 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2682
timestamp 1711653199
transform 1 0 2764 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1711653199
transform 1 0 2604 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1711653199
transform 1 0 2524 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1711653199
transform 1 0 2444 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2686
timestamp 1711653199
transform 1 0 2396 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1711653199
transform 1 0 1684 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_2688
timestamp 1711653199
transform 1 0 1676 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1711653199
transform 1 0 1636 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1711653199
transform 1 0 1604 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1711653199
transform 1 0 1508 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1711653199
transform 1 0 1492 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1711653199
transform 1 0 1772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2694
timestamp 1711653199
transform 1 0 1548 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1711653199
transform 1 0 2412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2696
timestamp 1711653199
transform 1 0 1556 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1711653199
transform 1 0 2780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2698
timestamp 1711653199
transform 1 0 2732 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2699
timestamp 1711653199
transform 1 0 2580 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1711653199
transform 1 0 2476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1711653199
transform 1 0 2420 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1711653199
transform 1 0 2404 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1711653199
transform 1 0 2436 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2704
timestamp 1711653199
transform 1 0 2436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1711653199
transform 1 0 2388 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1711653199
transform 1 0 1188 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1711653199
transform 1 0 2812 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2708
timestamp 1711653199
transform 1 0 2396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1711653199
transform 1 0 2492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2710
timestamp 1711653199
transform 1 0 2356 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1711653199
transform 1 0 2340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1711653199
transform 1 0 2284 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1711653199
transform 1 0 2228 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1711653199
transform 1 0 2164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1711653199
transform 1 0 2164 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1711653199
transform 1 0 2300 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2717
timestamp 1711653199
transform 1 0 2276 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1711653199
transform 1 0 2260 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1711653199
transform 1 0 2460 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1711653199
transform 1 0 2460 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1711653199
transform 1 0 2420 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1711653199
transform 1 0 2300 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1711653199
transform 1 0 3052 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1711653199
transform 1 0 2996 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1711653199
transform 1 0 2996 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1711653199
transform 1 0 2956 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1711653199
transform 1 0 2500 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1711653199
transform 1 0 2444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1711653199
transform 1 0 2500 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1711653199
transform 1 0 2300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2731
timestamp 1711653199
transform 1 0 2276 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1711653199
transform 1 0 2276 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2733
timestamp 1711653199
transform 1 0 2244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1711653199
transform 1 0 2204 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1711653199
transform 1 0 2172 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1711653199
transform 1 0 2164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1711653199
transform 1 0 2172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1711653199
transform 1 0 1876 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_2739
timestamp 1711653199
transform 1 0 2348 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1711653199
transform 1 0 2140 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1711653199
transform 1 0 2300 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1711653199
transform 1 0 2076 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1711653199
transform 1 0 2036 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2744
timestamp 1711653199
transform 1 0 1972 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1711653199
transform 1 0 1956 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2746
timestamp 1711653199
transform 1 0 2084 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1711653199
transform 1 0 1956 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1711653199
transform 1 0 1940 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1711653199
transform 1 0 2436 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1711653199
transform 1 0 2332 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1711653199
transform 1 0 2532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1711653199
transform 1 0 2420 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1711653199
transform 1 0 2468 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1711653199
transform 1 0 2468 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1711653199
transform 1 0 2420 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1711653199
transform 1 0 2532 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1711653199
transform 1 0 2452 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1711653199
transform 1 0 2412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1711653199
transform 1 0 2452 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1711653199
transform 1 0 2444 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1711653199
transform 1 0 2436 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1711653199
transform 1 0 3100 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2763
timestamp 1711653199
transform 1 0 2796 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2764
timestamp 1711653199
transform 1 0 2812 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1711653199
transform 1 0 2804 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1711653199
transform 1 0 2772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2767
timestamp 1711653199
transform 1 0 2772 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1711653199
transform 1 0 2756 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1711653199
transform 1 0 2756 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1711653199
transform 1 0 2828 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1711653199
transform 1 0 2812 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1711653199
transform 1 0 2804 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1711653199
transform 1 0 2804 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1711653199
transform 1 0 2796 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1711653199
transform 1 0 2596 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1711653199
transform 1 0 2580 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2777
timestamp 1711653199
transform 1 0 2564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1711653199
transform 1 0 2564 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2779
timestamp 1711653199
transform 1 0 2524 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1711653199
transform 1 0 2332 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2781
timestamp 1711653199
transform 1 0 3076 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1711653199
transform 1 0 3076 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1711653199
transform 1 0 3060 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1711653199
transform 1 0 3044 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2785
timestamp 1711653199
transform 1 0 2948 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2786
timestamp 1711653199
transform 1 0 2404 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2787
timestamp 1711653199
transform 1 0 1580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1711653199
transform 1 0 1564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1711653199
transform 1 0 3196 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2790
timestamp 1711653199
transform 1 0 3100 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1711653199
transform 1 0 3084 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1711653199
transform 1 0 3300 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1711653199
transform 1 0 3156 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2794
timestamp 1711653199
transform 1 0 3292 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2795
timestamp 1711653199
transform 1 0 3252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1711653199
transform 1 0 3228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1711653199
transform 1 0 3228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1711653199
transform 1 0 3316 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1711653199
transform 1 0 3316 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1711653199
transform 1 0 3268 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_2801
timestamp 1711653199
transform 1 0 1132 0 1 955
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1711653199
transform 1 0 612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1711653199
transform 1 0 1188 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1711653199
transform 1 0 1172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1711653199
transform 1 0 1164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1711653199
transform 1 0 1164 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1711653199
transform 1 0 1140 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2808
timestamp 1711653199
transform 1 0 1020 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1711653199
transform 1 0 3188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1711653199
transform 1 0 3172 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1711653199
transform 1 0 3012 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1711653199
transform 1 0 3012 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1711653199
transform 1 0 2980 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1711653199
transform 1 0 2972 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2815
timestamp 1711653199
transform 1 0 2660 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2816
timestamp 1711653199
transform 1 0 1724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1711653199
transform 1 0 1196 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1711653199
transform 1 0 1140 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2819
timestamp 1711653199
transform 1 0 1100 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2820
timestamp 1711653199
transform 1 0 1068 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1711653199
transform 1 0 1020 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1711653199
transform 1 0 980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1711653199
transform 1 0 1012 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1711653199
transform 1 0 972 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1711653199
transform 1 0 948 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2826
timestamp 1711653199
transform 1 0 876 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2827
timestamp 1711653199
transform 1 0 780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1711653199
transform 1 0 1060 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1711653199
transform 1 0 1060 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2830
timestamp 1711653199
transform 1 0 1020 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1711653199
transform 1 0 1012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1711653199
transform 1 0 1132 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2833
timestamp 1711653199
transform 1 0 300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2834
timestamp 1711653199
transform 1 0 1244 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1711653199
transform 1 0 1220 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2836
timestamp 1711653199
transform 1 0 1268 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1711653199
transform 1 0 1220 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1711653199
transform 1 0 1324 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2839
timestamp 1711653199
transform 1 0 1316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1711653199
transform 1 0 252 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1711653199
transform 1 0 228 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2842
timestamp 1711653199
transform 1 0 212 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2843
timestamp 1711653199
transform 1 0 420 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_2844
timestamp 1711653199
transform 1 0 332 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_2845
timestamp 1711653199
transform 1 0 316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2846
timestamp 1711653199
transform 1 0 532 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1711653199
transform 1 0 308 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1711653199
transform 1 0 644 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2849
timestamp 1711653199
transform 1 0 572 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2850
timestamp 1711653199
transform 1 0 2532 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2851
timestamp 1711653199
transform 1 0 2508 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2852
timestamp 1711653199
transform 1 0 700 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1711653199
transform 1 0 596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1711653199
transform 1 0 516 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1711653199
transform 1 0 724 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1711653199
transform 1 0 668 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1711653199
transform 1 0 692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1711653199
transform 1 0 692 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1711653199
transform 1 0 644 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1711653199
transform 1 0 644 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1711653199
transform 1 0 812 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1711653199
transform 1 0 740 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1711653199
transform 1 0 628 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1711653199
transform 1 0 308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2865
timestamp 1711653199
transform 1 0 276 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1711653199
transform 1 0 348 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1711653199
transform 1 0 324 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1711653199
transform 1 0 380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_2869
timestamp 1711653199
transform 1 0 332 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2870
timestamp 1711653199
transform 1 0 156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2871
timestamp 1711653199
transform 1 0 444 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2872
timestamp 1711653199
transform 1 0 388 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2873
timestamp 1711653199
transform 1 0 276 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2874
timestamp 1711653199
transform 1 0 148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1711653199
transform 1 0 324 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2876
timestamp 1711653199
transform 1 0 252 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1711653199
transform 1 0 220 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1711653199
transform 1 0 2396 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1711653199
transform 1 0 2396 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1711653199
transform 1 0 2484 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1711653199
transform 1 0 2388 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1711653199
transform 1 0 2508 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1711653199
transform 1 0 2412 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_2884
timestamp 1711653199
transform 1 0 2548 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2885
timestamp 1711653199
transform 1 0 2540 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1711653199
transform 1 0 2652 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1711653199
transform 1 0 2556 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1711653199
transform 1 0 2652 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1711653199
transform 1 0 620 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2890
timestamp 1711653199
transform 1 0 532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1711653199
transform 1 0 356 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2892
timestamp 1711653199
transform 1 0 588 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1711653199
transform 1 0 556 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1711653199
transform 1 0 644 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1711653199
transform 1 0 620 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1711653199
transform 1 0 732 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2897
timestamp 1711653199
transform 1 0 660 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1711653199
transform 1 0 628 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1711653199
transform 1 0 668 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1711653199
transform 1 0 660 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_2901
timestamp 1711653199
transform 1 0 548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1711653199
transform 1 0 540 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1711653199
transform 1 0 516 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1711653199
transform 1 0 460 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2905
timestamp 1711653199
transform 1 0 356 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1711653199
transform 1 0 300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2907
timestamp 1711653199
transform 1 0 412 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2908
timestamp 1711653199
transform 1 0 388 0 1 685
box -2 -2 2 2
use M2_M1  M2_M1_2909
timestamp 1711653199
transform 1 0 380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2910
timestamp 1711653199
transform 1 0 324 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1711653199
transform 1 0 284 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_2912
timestamp 1711653199
transform 1 0 524 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2913
timestamp 1711653199
transform 1 0 428 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2914
timestamp 1711653199
transform 1 0 380 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2915
timestamp 1711653199
transform 1 0 284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1711653199
transform 1 0 132 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2917
timestamp 1711653199
transform 1 0 132 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1711653199
transform 1 0 116 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1711653199
transform 1 0 116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2920
timestamp 1711653199
transform 1 0 324 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1711653199
transform 1 0 324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2922
timestamp 1711653199
transform 1 0 284 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1711653199
transform 1 0 2860 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1711653199
transform 1 0 2660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2925
timestamp 1711653199
transform 1 0 2612 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1711653199
transform 1 0 2740 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2927
timestamp 1711653199
transform 1 0 2532 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1711653199
transform 1 0 2500 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_2929
timestamp 1711653199
transform 1 0 1068 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2930
timestamp 1711653199
transform 1 0 972 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2931
timestamp 1711653199
transform 1 0 948 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2932
timestamp 1711653199
transform 1 0 1052 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1711653199
transform 1 0 1036 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2934
timestamp 1711653199
transform 1 0 1052 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1711653199
transform 1 0 1036 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1711653199
transform 1 0 980 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_2937
timestamp 1711653199
transform 1 0 908 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2938
timestamp 1711653199
transform 1 0 908 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1711653199
transform 1 0 1076 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1711653199
transform 1 0 1076 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2941
timestamp 1711653199
transform 1 0 1044 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1711653199
transform 1 0 1276 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1711653199
transform 1 0 1092 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1711653199
transform 1 0 1060 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1711653199
transform 1 0 868 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1711653199
transform 1 0 284 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2947
timestamp 1711653199
transform 1 0 1252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2948
timestamp 1711653199
transform 1 0 956 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2949
timestamp 1711653199
transform 1 0 1356 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1711653199
transform 1 0 1196 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1711653199
transform 1 0 1196 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1711653199
transform 1 0 1292 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1711653199
transform 1 0 1268 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1711653199
transform 1 0 1268 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2955
timestamp 1711653199
transform 1 0 212 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1711653199
transform 1 0 212 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1711653199
transform 1 0 180 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1711653199
transform 1 0 460 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1711653199
transform 1 0 364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1711653199
transform 1 0 332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1711653199
transform 1 0 2972 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1711653199
transform 1 0 2796 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1711653199
transform 1 0 3308 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1711653199
transform 1 0 2972 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1711653199
transform 1 0 3380 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1711653199
transform 1 0 3380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1711653199
transform 1 0 3324 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1711653199
transform 1 0 3292 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1711653199
transform 1 0 3380 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1711653199
transform 1 0 3340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1711653199
transform 1 0 3340 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1711653199
transform 1 0 3116 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1711653199
transform 1 0 3004 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1711653199
transform 1 0 2980 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2975
timestamp 1711653199
transform 1 0 2468 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1711653199
transform 1 0 2332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1711653199
transform 1 0 2268 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1711653199
transform 1 0 2260 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2979
timestamp 1711653199
transform 1 0 2236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1711653199
transform 1 0 2076 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1711653199
transform 1 0 2660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1711653199
transform 1 0 2564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2983
timestamp 1711653199
transform 1 0 2532 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1711653199
transform 1 0 2468 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1711653199
transform 1 0 2396 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1711653199
transform 1 0 2324 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2987
timestamp 1711653199
transform 1 0 2260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1711653199
transform 1 0 1900 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1711653199
transform 1 0 1484 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1711653199
transform 1 0 1484 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1711653199
transform 1 0 1484 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1711653199
transform 1 0 2100 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1711653199
transform 1 0 2036 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1711653199
transform 1 0 1964 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1711653199
transform 1 0 2084 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1711653199
transform 1 0 1852 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1711653199
transform 1 0 1748 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1711653199
transform 1 0 2228 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1711653199
transform 1 0 1924 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1711653199
transform 1 0 1892 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1711653199
transform 1 0 2340 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1711653199
transform 1 0 2324 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1711653199
transform 1 0 2308 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1711653199
transform 1 0 2276 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1711653199
transform 1 0 2244 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3006
timestamp 1711653199
transform 1 0 2436 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1711653199
transform 1 0 2428 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1711653199
transform 1 0 2300 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1711653199
transform 1 0 2500 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1711653199
transform 1 0 2196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3011
timestamp 1711653199
transform 1 0 2196 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1711653199
transform 1 0 2324 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1711653199
transform 1 0 2132 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1711653199
transform 1 0 2132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3015
timestamp 1711653199
transform 1 0 2516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3016
timestamp 1711653199
transform 1 0 2356 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1711653199
transform 1 0 2356 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3018
timestamp 1711653199
transform 1 0 1772 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1711653199
transform 1 0 1684 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1711653199
transform 1 0 1820 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1711653199
transform 1 0 1724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1711653199
transform 1 0 1924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1711653199
transform 1 0 1844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1711653199
transform 1 0 2556 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1711653199
transform 1 0 1900 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3026
timestamp 1711653199
transform 1 0 2868 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1711653199
transform 1 0 2820 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1711653199
transform 1 0 2804 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1711653199
transform 1 0 2540 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1711653199
transform 1 0 2684 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1711653199
transform 1 0 2684 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1711653199
transform 1 0 2644 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1711653199
transform 1 0 2548 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1711653199
transform 1 0 2628 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1711653199
transform 1 0 2572 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1711653199
transform 1 0 2524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1711653199
transform 1 0 1868 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1711653199
transform 1 0 1660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1711653199
transform 1 0 1532 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3040
timestamp 1711653199
transform 1 0 1956 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3041
timestamp 1711653199
transform 1 0 1892 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1711653199
transform 1 0 1636 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1711653199
transform 1 0 2036 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1711653199
transform 1 0 1740 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1711653199
transform 1 0 1748 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1711653199
transform 1 0 788 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1711653199
transform 1 0 1796 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1711653199
transform 1 0 1748 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1711653199
transform 1 0 1724 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1711653199
transform 1 0 1196 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3051
timestamp 1711653199
transform 1 0 2804 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1711653199
transform 1 0 1780 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1711653199
transform 1 0 3084 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1711653199
transform 1 0 2780 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3055
timestamp 1711653199
transform 1 0 2956 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1711653199
transform 1 0 2876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1711653199
transform 1 0 2844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3058
timestamp 1711653199
transform 1 0 2700 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1711653199
transform 1 0 2508 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1711653199
transform 1 0 2468 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3061
timestamp 1711653199
transform 1 0 2452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3062
timestamp 1711653199
transform 1 0 2444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1711653199
transform 1 0 3212 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1711653199
transform 1 0 3084 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3065
timestamp 1711653199
transform 1 0 3036 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1711653199
transform 1 0 3356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1711653199
transform 1 0 3340 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1711653199
transform 1 0 3332 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1711653199
transform 1 0 3316 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1711653199
transform 1 0 3228 0 1 1255
box -2 -2 2 2
use M2_M1  M2_M1_3071
timestamp 1711653199
transform 1 0 3396 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_3072
timestamp 1711653199
transform 1 0 3364 0 1 1203
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1711653199
transform 1 0 3236 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1711653199
transform 1 0 1124 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1711653199
transform 1 0 308 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1711653199
transform 1 0 1244 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1711653199
transform 1 0 1148 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1711653199
transform 1 0 1172 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1711653199
transform 1 0 1092 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1711653199
transform 1 0 1060 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1711653199
transform 1 0 996 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1711653199
transform 1 0 940 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3083
timestamp 1711653199
transform 1 0 900 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1711653199
transform 1 0 876 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1711653199
transform 1 0 1124 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1711653199
transform 1 0 1004 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1711653199
transform 1 0 860 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1711653199
transform 1 0 892 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1711653199
transform 1 0 780 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1711653199
transform 1 0 772 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1711653199
transform 1 0 1412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3092
timestamp 1711653199
transform 1 0 1380 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1711653199
transform 1 0 1220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3094
timestamp 1711653199
transform 1 0 1260 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1711653199
transform 1 0 1188 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1711653199
transform 1 0 1188 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1711653199
transform 1 0 324 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1711653199
transform 1 0 284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1711653199
transform 1 0 284 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3100
timestamp 1711653199
transform 1 0 428 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1711653199
transform 1 0 332 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1711653199
transform 1 0 740 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1711653199
transform 1 0 388 0 1 1445
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1711653199
transform 1 0 780 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1711653199
transform 1 0 748 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1711653199
transform 1 0 796 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1711653199
transform 1 0 772 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1711653199
transform 1 0 732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1711653199
transform 1 0 628 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1711653199
transform 1 0 612 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1711653199
transform 1 0 980 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1711653199
transform 1 0 788 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1711653199
transform 1 0 692 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1711653199
transform 1 0 684 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3115
timestamp 1711653199
transform 1 0 612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1711653199
transform 1 0 380 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1711653199
transform 1 0 204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1711653199
transform 1 0 444 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1711653199
transform 1 0 420 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1711653199
transform 1 0 476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1711653199
transform 1 0 420 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1711653199
transform 1 0 348 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1711653199
transform 1 0 580 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1711653199
transform 1 0 484 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3125
timestamp 1711653199
transform 1 0 172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1711653199
transform 1 0 164 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1711653199
transform 1 0 164 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3128
timestamp 1711653199
transform 1 0 220 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1711653199
transform 1 0 220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3130
timestamp 1711653199
transform 1 0 196 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3131
timestamp 1711653199
transform 1 0 196 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1711653199
transform 1 0 2036 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3133
timestamp 1711653199
transform 1 0 2004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3134
timestamp 1711653199
transform 1 0 2012 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3135
timestamp 1711653199
transform 1 0 1852 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3136
timestamp 1711653199
transform 1 0 1852 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1711653199
transform 1 0 1844 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3138
timestamp 1711653199
transform 1 0 2108 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3139
timestamp 1711653199
transform 1 0 2004 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3140
timestamp 1711653199
transform 1 0 1820 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3141
timestamp 1711653199
transform 1 0 1860 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3142
timestamp 1711653199
transform 1 0 1724 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1711653199
transform 1 0 1628 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1711653199
transform 1 0 1836 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1711653199
transform 1 0 1836 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3146
timestamp 1711653199
transform 1 0 1804 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1711653199
transform 1 0 1796 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3148
timestamp 1711653199
transform 1 0 2188 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1711653199
transform 1 0 2036 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1711653199
transform 1 0 2060 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1711653199
transform 1 0 2012 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3152
timestamp 1711653199
transform 1 0 2116 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1711653199
transform 1 0 1956 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1711653199
transform 1 0 1908 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3155
timestamp 1711653199
transform 1 0 2028 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1711653199
transform 1 0 1668 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1711653199
transform 1 0 2332 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3158
timestamp 1711653199
transform 1 0 2228 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3159
timestamp 1711653199
transform 1 0 2172 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1711653199
transform 1 0 2284 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1711653199
transform 1 0 2204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1711653199
transform 1 0 2204 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1711653199
transform 1 0 1484 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1711653199
transform 1 0 1452 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1711653199
transform 1 0 1444 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1711653199
transform 1 0 1444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1711653199
transform 1 0 1724 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1711653199
transform 1 0 1412 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1711653199
transform 1 0 1452 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1711653199
transform 1 0 1412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1711653199
transform 1 0 1428 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3172
timestamp 1711653199
transform 1 0 1124 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1711653199
transform 1 0 1116 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1711653199
transform 1 0 996 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1711653199
transform 1 0 2308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1711653199
transform 1 0 2292 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1711653199
transform 1 0 2292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1711653199
transform 1 0 2228 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1711653199
transform 1 0 1532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1711653199
transform 1 0 948 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3181
timestamp 1711653199
transform 1 0 900 0 1 1045
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1711653199
transform 1 0 900 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1711653199
transform 1 0 900 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3184
timestamp 1711653199
transform 1 0 1364 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1711653199
transform 1 0 1308 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3186
timestamp 1711653199
transform 1 0 980 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3187
timestamp 1711653199
transform 1 0 972 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1711653199
transform 1 0 972 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3189
timestamp 1711653199
transform 1 0 956 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1711653199
transform 1 0 1028 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1711653199
transform 1 0 1004 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3192
timestamp 1711653199
transform 1 0 948 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1711653199
transform 1 0 668 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3194
timestamp 1711653199
transform 1 0 668 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1711653199
transform 1 0 628 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1711653199
transform 1 0 1348 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1711653199
transform 1 0 1228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1711653199
transform 1 0 3204 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1711653199
transform 1 0 3076 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1711653199
transform 1 0 2956 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1711653199
transform 1 0 2756 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1711653199
transform 1 0 2716 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3203
timestamp 1711653199
transform 1 0 1300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1711653199
transform 1 0 1228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1711653199
transform 1 0 1188 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1711653199
transform 1 0 1444 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1711653199
transform 1 0 1324 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3208
timestamp 1711653199
transform 1 0 1252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1711653199
transform 1 0 1244 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3210
timestamp 1711653199
transform 1 0 1212 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1711653199
transform 1 0 1196 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1711653199
transform 1 0 1492 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1711653199
transform 1 0 1388 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3214
timestamp 1711653199
transform 1 0 1284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1711653199
transform 1 0 1276 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1711653199
transform 1 0 1244 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1711653199
transform 1 0 1180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1711653199
transform 1 0 860 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1711653199
transform 1 0 820 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1711653199
transform 1 0 804 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1711653199
transform 1 0 1244 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1711653199
transform 1 0 836 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1711653199
transform 1 0 836 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1711653199
transform 1 0 636 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3225
timestamp 1711653199
transform 1 0 556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3226
timestamp 1711653199
transform 1 0 524 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3227
timestamp 1711653199
transform 1 0 1820 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1711653199
transform 1 0 1724 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1711653199
transform 1 0 2036 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1711653199
transform 1 0 1796 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1711653199
transform 1 0 2044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1711653199
transform 1 0 1956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3233
timestamp 1711653199
transform 1 0 1972 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3234
timestamp 1711653199
transform 1 0 1940 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1711653199
transform 1 0 1940 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1711653199
transform 1 0 1932 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3237
timestamp 1711653199
transform 1 0 1836 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1711653199
transform 1 0 1812 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1711653199
transform 1 0 1948 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1711653199
transform 1 0 1948 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1711653199
transform 1 0 1948 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1711653199
transform 1 0 1892 0 1 1655
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1711653199
transform 1 0 1892 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1711653199
transform 1 0 1892 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_3245
timestamp 1711653199
transform 1 0 1868 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1711653199
transform 1 0 1868 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1711653199
transform 1 0 1164 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1711653199
transform 1 0 1140 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1711653199
transform 1 0 2236 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1711653199
transform 1 0 2108 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1711653199
transform 1 0 2100 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1711653199
transform 1 0 2036 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1711653199
transform 1 0 1996 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1711653199
transform 1 0 1628 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1711653199
transform 1 0 812 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1711653199
transform 1 0 1988 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1711653199
transform 1 0 1884 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1711653199
transform 1 0 1876 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1711653199
transform 1 0 1836 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1711653199
transform 1 0 1700 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1711653199
transform 1 0 1644 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1711653199
transform 1 0 1876 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1711653199
transform 1 0 1860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1711653199
transform 1 0 1868 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1711653199
transform 1 0 1036 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1711653199
transform 1 0 876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1711653199
transform 1 0 676 0 1 1445
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1711653199
transform 1 0 564 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1711653199
transform 1 0 524 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1711653199
transform 1 0 2964 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1711653199
transform 1 0 2956 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1711653199
transform 1 0 2932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1711653199
transform 1 0 2908 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1711653199
transform 1 0 2844 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1711653199
transform 1 0 1988 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1711653199
transform 1 0 1892 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3277
timestamp 1711653199
transform 1 0 1892 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1711653199
transform 1 0 2556 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1711653199
transform 1 0 2516 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1711653199
transform 1 0 2300 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1711653199
transform 1 0 2228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3282
timestamp 1711653199
transform 1 0 2084 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1711653199
transform 1 0 1932 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1711653199
transform 1 0 1764 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1711653199
transform 1 0 1732 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1711653199
transform 1 0 1732 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1711653199
transform 1 0 1732 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1711653199
transform 1 0 1692 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1711653199
transform 1 0 1388 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1711653199
transform 1 0 1076 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1711653199
transform 1 0 1524 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1711653199
transform 1 0 1412 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1711653199
transform 1 0 1452 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1711653199
transform 1 0 1428 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3295
timestamp 1711653199
transform 1 0 1668 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1711653199
transform 1 0 1380 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1711653199
transform 1 0 1404 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1711653199
transform 1 0 292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3299
timestamp 1711653199
transform 1 0 252 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3300
timestamp 1711653199
transform 1 0 212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1711653199
transform 1 0 196 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1711653199
transform 1 0 172 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1711653199
transform 1 0 308 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3304
timestamp 1711653199
transform 1 0 284 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1711653199
transform 1 0 476 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1711653199
transform 1 0 468 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3307
timestamp 1711653199
transform 1 0 420 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1711653199
transform 1 0 412 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1711653199
transform 1 0 364 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1711653199
transform 1 0 300 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1711653199
transform 1 0 1340 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3312
timestamp 1711653199
transform 1 0 1316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1711653199
transform 1 0 332 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1711653199
transform 1 0 124 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1711653199
transform 1 0 124 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3316
timestamp 1711653199
transform 1 0 636 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1711653199
transform 1 0 332 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1711653199
transform 1 0 332 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1711653199
transform 1 0 324 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1711653199
transform 1 0 316 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3321
timestamp 1711653199
transform 1 0 308 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1711653199
transform 1 0 300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1711653199
transform 1 0 236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1711653199
transform 1 0 1660 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3325
timestamp 1711653199
transform 1 0 1652 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1711653199
transform 1 0 2244 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1711653199
transform 1 0 1724 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1711653199
transform 1 0 2228 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3329
timestamp 1711653199
transform 1 0 2228 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1711653199
transform 1 0 2868 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1711653199
transform 1 0 2604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1711653199
transform 1 0 2580 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1711653199
transform 1 0 2324 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1711653199
transform 1 0 2180 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1711653199
transform 1 0 1444 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1711653199
transform 1 0 1428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1711653199
transform 1 0 2244 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1711653199
transform 1 0 2244 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3339
timestamp 1711653199
transform 1 0 2212 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3340
timestamp 1711653199
transform 1 0 2148 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1711653199
transform 1 0 2124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1711653199
transform 1 0 1940 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1711653199
transform 1 0 1940 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1711653199
transform 1 0 1932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1711653199
transform 1 0 2252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1711653199
transform 1 0 2196 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1711653199
transform 1 0 2172 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1711653199
transform 1 0 2108 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3349
timestamp 1711653199
transform 1 0 2044 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1711653199
transform 1 0 3060 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1711653199
transform 1 0 1644 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3352
timestamp 1711653199
transform 1 0 2748 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3353
timestamp 1711653199
transform 1 0 2700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1711653199
transform 1 0 2684 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1711653199
transform 1 0 1684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1711653199
transform 1 0 1668 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3357
timestamp 1711653199
transform 1 0 1628 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1711653199
transform 1 0 1684 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1711653199
transform 1 0 1484 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1711653199
transform 1 0 1484 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1711653199
transform 1 0 1436 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1711653199
transform 1 0 1436 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1711653199
transform 1 0 1420 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1711653199
transform 1 0 1412 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_3365
timestamp 1711653199
transform 1 0 3044 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1711653199
transform 1 0 3028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3367
timestamp 1711653199
transform 1 0 3028 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1711653199
transform 1 0 2956 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1711653199
transform 1 0 2916 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3370
timestamp 1711653199
transform 1 0 2916 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1711653199
transform 1 0 2436 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1711653199
transform 1 0 2372 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1711653199
transform 1 0 3124 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1711653199
transform 1 0 3084 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1711653199
transform 1 0 3348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3376
timestamp 1711653199
transform 1 0 3276 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1711653199
transform 1 0 3252 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3378
timestamp 1711653199
transform 1 0 3244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1711653199
transform 1 0 3116 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1711653199
transform 1 0 2860 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1711653199
transform 1 0 3284 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1711653199
transform 1 0 3236 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1711653199
transform 1 0 3236 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1711653199
transform 1 0 3236 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1711653199
transform 1 0 3140 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3386
timestamp 1711653199
transform 1 0 2988 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3387
timestamp 1711653199
transform 1 0 1524 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3388
timestamp 1711653199
transform 1 0 1492 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1711653199
transform 1 0 1508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1711653199
transform 1 0 1484 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1711653199
transform 1 0 1484 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1711653199
transform 1 0 1172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1711653199
transform 1 0 2868 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1711653199
transform 1 0 2868 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1711653199
transform 1 0 2852 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1711653199
transform 1 0 2780 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1711653199
transform 1 0 2764 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1711653199
transform 1 0 2764 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1711653199
transform 1 0 1100 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1711653199
transform 1 0 1052 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1711653199
transform 1 0 916 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3402
timestamp 1711653199
transform 1 0 1372 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1711653199
transform 1 0 1164 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1711653199
transform 1 0 1164 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1711653199
transform 1 0 1164 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1711653199
transform 1 0 1124 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1711653199
transform 1 0 1124 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1711653199
transform 1 0 1076 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3409
timestamp 1711653199
transform 1 0 1452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3410
timestamp 1711653199
transform 1 0 1436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1711653199
transform 1 0 1188 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1711653199
transform 1 0 1140 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1711653199
transform 1 0 1108 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1711653199
transform 1 0 1068 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3415
timestamp 1711653199
transform 1 0 1180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3416
timestamp 1711653199
transform 1 0 1044 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3417
timestamp 1711653199
transform 1 0 916 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1711653199
transform 1 0 892 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_3419
timestamp 1711653199
transform 1 0 732 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3420
timestamp 1711653199
transform 1 0 588 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_3421
timestamp 1711653199
transform 1 0 1508 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_3422
timestamp 1711653199
transform 1 0 540 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3423
timestamp 1711653199
transform 1 0 1340 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3424
timestamp 1711653199
transform 1 0 932 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3425
timestamp 1711653199
transform 1 0 540 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_3426
timestamp 1711653199
transform 1 0 540 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_3427
timestamp 1711653199
transform 1 0 532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1711653199
transform 1 0 524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3429
timestamp 1711653199
transform 1 0 524 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3430
timestamp 1711653199
transform 1 0 468 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1711653199
transform 1 0 740 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1711653199
transform 1 0 516 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1711653199
transform 1 0 516 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3434
timestamp 1711653199
transform 1 0 500 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3435
timestamp 1711653199
transform 1 0 388 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3436
timestamp 1711653199
transform 1 0 380 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1711653199
transform 1 0 372 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3438
timestamp 1711653199
transform 1 0 1428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1711653199
transform 1 0 876 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1711653199
transform 1 0 772 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_3441
timestamp 1711653199
transform 1 0 580 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3442
timestamp 1711653199
transform 1 0 564 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3443
timestamp 1711653199
transform 1 0 516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1711653199
transform 1 0 572 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1711653199
transform 1 0 548 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3446
timestamp 1711653199
transform 1 0 340 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1711653199
transform 1 0 260 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1711653199
transform 1 0 252 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_3449
timestamp 1711653199
transform 1 0 236 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1711653199
transform 1 0 1580 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1711653199
transform 1 0 1540 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3452
timestamp 1711653199
transform 1 0 1652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1711653199
transform 1 0 1628 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1711653199
transform 1 0 1668 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3455
timestamp 1711653199
transform 1 0 1588 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1711653199
transform 1 0 2396 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1711653199
transform 1 0 1732 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1711653199
transform 1 0 2348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1711653199
transform 1 0 2348 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1711653199
transform 1 0 2460 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3461
timestamp 1711653199
transform 1 0 2380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3462
timestamp 1711653199
transform 1 0 2668 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1711653199
transform 1 0 2388 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1711653199
transform 1 0 2676 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1711653199
transform 1 0 2676 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1711653199
transform 1 0 2684 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3467
timestamp 1711653199
transform 1 0 788 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3468
timestamp 1711653199
transform 1 0 716 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3469
timestamp 1711653199
transform 1 0 388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1711653199
transform 1 0 708 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3471
timestamp 1711653199
transform 1 0 708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3472
timestamp 1711653199
transform 1 0 700 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3473
timestamp 1711653199
transform 1 0 636 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1711653199
transform 1 0 620 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3475
timestamp 1711653199
transform 1 0 612 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1711653199
transform 1 0 612 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1711653199
transform 1 0 676 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3478
timestamp 1711653199
transform 1 0 668 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1711653199
transform 1 0 620 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1711653199
transform 1 0 324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3481
timestamp 1711653199
transform 1 0 308 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1711653199
transform 1 0 404 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3483
timestamp 1711653199
transform 1 0 404 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1711653199
transform 1 0 484 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1711653199
transform 1 0 332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3486
timestamp 1711653199
transform 1 0 228 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3487
timestamp 1711653199
transform 1 0 460 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1711653199
transform 1 0 460 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1711653199
transform 1 0 404 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3490
timestamp 1711653199
transform 1 0 260 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3491
timestamp 1711653199
transform 1 0 188 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3492
timestamp 1711653199
transform 1 0 132 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3493
timestamp 1711653199
transform 1 0 340 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3494
timestamp 1711653199
transform 1 0 252 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3495
timestamp 1711653199
transform 1 0 180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3496
timestamp 1711653199
transform 1 0 2572 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3497
timestamp 1711653199
transform 1 0 2492 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3498
timestamp 1711653199
transform 1 0 2820 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1711653199
transform 1 0 2604 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3500
timestamp 1711653199
transform 1 0 2556 0 1 105
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1711653199
transform 1 0 1148 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1711653199
transform 1 0 1052 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3503
timestamp 1711653199
transform 1 0 1028 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3504
timestamp 1711653199
transform 1 0 1124 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3505
timestamp 1711653199
transform 1 0 1084 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1711653199
transform 1 0 1108 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3507
timestamp 1711653199
transform 1 0 956 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3508
timestamp 1711653199
transform 1 0 916 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1711653199
transform 1 0 764 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3510
timestamp 1711653199
transform 1 0 756 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3511
timestamp 1711653199
transform 1 0 996 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3512
timestamp 1711653199
transform 1 0 972 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1711653199
transform 1 0 932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3514
timestamp 1711653199
transform 1 0 940 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1711653199
transform 1 0 364 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1711653199
transform 1 0 1172 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3517
timestamp 1711653199
transform 1 0 1020 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1711653199
transform 1 0 1276 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3519
timestamp 1711653199
transform 1 0 1276 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3520
timestamp 1711653199
transform 1 0 1156 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1711653199
transform 1 0 1188 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1711653199
transform 1 0 1188 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1711653199
transform 1 0 340 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1711653199
transform 1 0 276 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3525
timestamp 1711653199
transform 1 0 188 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3526
timestamp 1711653199
transform 1 0 420 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1711653199
transform 1 0 404 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1711653199
transform 1 0 3100 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3529
timestamp 1711653199
transform 1 0 2860 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3530
timestamp 1711653199
transform 1 0 3188 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1711653199
transform 1 0 3164 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3532
timestamp 1711653199
transform 1 0 3180 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3533
timestamp 1711653199
transform 1 0 3172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1711653199
transform 1 0 3172 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3535
timestamp 1711653199
transform 1 0 3380 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1711653199
transform 1 0 3220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3537
timestamp 1711653199
transform 1 0 3204 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1711653199
transform 1 0 3068 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3539
timestamp 1711653199
transform 1 0 3060 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3540
timestamp 1711653199
transform 1 0 2996 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1711653199
transform 1 0 2972 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3542
timestamp 1711653199
transform 1 0 2540 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3543
timestamp 1711653199
transform 1 0 2468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3544
timestamp 1711653199
transform 1 0 2436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1711653199
transform 1 0 2220 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1711653199
transform 1 0 2780 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1711653199
transform 1 0 2628 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1711653199
transform 1 0 2564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3549
timestamp 1711653199
transform 1 0 2524 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1711653199
transform 1 0 2780 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1711653199
transform 1 0 2660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3552
timestamp 1711653199
transform 1 0 2652 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1711653199
transform 1 0 2596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1711653199
transform 1 0 2588 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1711653199
transform 1 0 2548 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3556
timestamp 1711653199
transform 1 0 2356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3557
timestamp 1711653199
transform 1 0 2356 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1711653199
transform 1 0 2444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1711653199
transform 1 0 2444 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1711653199
transform 1 0 2340 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1711653199
transform 1 0 2476 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3562
timestamp 1711653199
transform 1 0 2164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3563
timestamp 1711653199
transform 1 0 2292 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3564
timestamp 1711653199
transform 1 0 2188 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3565
timestamp 1711653199
transform 1 0 2164 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1711653199
transform 1 0 2500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3567
timestamp 1711653199
transform 1 0 2492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3568
timestamp 1711653199
transform 1 0 2436 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3569
timestamp 1711653199
transform 1 0 2404 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3570
timestamp 1711653199
transform 1 0 2396 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3571
timestamp 1711653199
transform 1 0 2516 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1711653199
transform 1 0 2516 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1711653199
transform 1 0 2500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3574
timestamp 1711653199
transform 1 0 2492 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3575
timestamp 1711653199
transform 1 0 2460 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1711653199
transform 1 0 2404 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1711653199
transform 1 0 2540 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1711653199
transform 1 0 2524 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1711653199
transform 1 0 1852 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3580
timestamp 1711653199
transform 1 0 1836 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1711653199
transform 1 0 1788 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3582
timestamp 1711653199
transform 1 0 1428 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1711653199
transform 1 0 940 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1711653199
transform 1 0 1748 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1711653199
transform 1 0 1652 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1711653199
transform 1 0 1652 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3587
timestamp 1711653199
transform 1 0 1388 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1711653199
transform 1 0 1588 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1711653199
transform 1 0 1588 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_3590
timestamp 1711653199
transform 1 0 1588 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1711653199
transform 1 0 1532 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3592
timestamp 1711653199
transform 1 0 1548 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1711653199
transform 1 0 1524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1711653199
transform 1 0 1508 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1711653199
transform 1 0 1468 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_3596
timestamp 1711653199
transform 1 0 1428 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1711653199
transform 1 0 1428 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1711653199
transform 1 0 1812 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1711653199
transform 1 0 1812 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3600
timestamp 1711653199
transform 1 0 1532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3601
timestamp 1711653199
transform 1 0 1388 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1711653199
transform 1 0 1404 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_3603
timestamp 1711653199
transform 1 0 1100 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1711653199
transform 1 0 1508 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_3605
timestamp 1711653199
transform 1 0 540 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1711653199
transform 1 0 500 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1711653199
transform 1 0 388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3608
timestamp 1711653199
transform 1 0 548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3609
timestamp 1711653199
transform 1 0 244 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1711653199
transform 1 0 244 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1711653199
transform 1 0 2068 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3612
timestamp 1711653199
transform 1 0 2060 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_3613
timestamp 1711653199
transform 1 0 1980 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1711653199
transform 1 0 1740 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1711653199
transform 1 0 1612 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1711653199
transform 1 0 1532 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_3617
timestamp 1711653199
transform 1 0 2236 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3618
timestamp 1711653199
transform 1 0 1548 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3619
timestamp 1711653199
transform 1 0 1500 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1711653199
transform 1 0 140 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3621
timestamp 1711653199
transform 1 0 1276 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3622
timestamp 1711653199
transform 1 0 212 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1711653199
transform 1 0 148 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3624
timestamp 1711653199
transform 1 0 124 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3625
timestamp 1711653199
transform 1 0 100 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3626
timestamp 1711653199
transform 1 0 172 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3627
timestamp 1711653199
transform 1 0 92 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1711653199
transform 1 0 84 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1711653199
transform 1 0 140 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1711653199
transform 1 0 92 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1711653199
transform 1 0 228 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3632
timestamp 1711653199
transform 1 0 172 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1711653199
transform 1 0 124 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3634
timestamp 1711653199
transform 1 0 324 0 1 1235
box -2 -2 2 2
use M2_M1  M2_M1_3635
timestamp 1711653199
transform 1 0 172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_3636
timestamp 1711653199
transform 1 0 164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_3637
timestamp 1711653199
transform 1 0 2364 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3638
timestamp 1711653199
transform 1 0 2212 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1711653199
transform 1 0 2364 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1711653199
transform 1 0 2284 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3641
timestamp 1711653199
transform 1 0 2460 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3642
timestamp 1711653199
transform 1 0 2356 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1711653199
transform 1 0 2292 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1711653199
transform 1 0 2292 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3645
timestamp 1711653199
transform 1 0 2412 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1711653199
transform 1 0 2380 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3647
timestamp 1711653199
transform 1 0 2324 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3648
timestamp 1711653199
transform 1 0 2260 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3649
timestamp 1711653199
transform 1 0 3084 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3650
timestamp 1711653199
transform 1 0 1604 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3651
timestamp 1711653199
transform 1 0 1628 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3652
timestamp 1711653199
transform 1 0 1380 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3653
timestamp 1711653199
transform 1 0 1260 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_3654
timestamp 1711653199
transform 1 0 3148 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3655
timestamp 1711653199
transform 1 0 3108 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3656
timestamp 1711653199
transform 1 0 3052 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3657
timestamp 1711653199
transform 1 0 3220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3658
timestamp 1711653199
transform 1 0 3116 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3659
timestamp 1711653199
transform 1 0 3356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3660
timestamp 1711653199
transform 1 0 3268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3661
timestamp 1711653199
transform 1 0 3212 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3662
timestamp 1711653199
transform 1 0 3364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3663
timestamp 1711653199
transform 1 0 3292 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3664
timestamp 1711653199
transform 1 0 3252 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3665
timestamp 1711653199
transform 1 0 1372 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1711653199
transform 1 0 1340 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3667
timestamp 1711653199
transform 1 0 1364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3668
timestamp 1711653199
transform 1 0 1060 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3669
timestamp 1711653199
transform 1 0 964 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3670
timestamp 1711653199
transform 1 0 860 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3671
timestamp 1711653199
transform 1 0 860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3672
timestamp 1711653199
transform 1 0 1020 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3673
timestamp 1711653199
transform 1 0 932 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3674
timestamp 1711653199
transform 1 0 1932 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_3675
timestamp 1711653199
transform 1 0 1932 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1711653199
transform 1 0 1588 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_3677
timestamp 1711653199
transform 1 0 1348 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3678
timestamp 1711653199
transform 1 0 1364 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3679
timestamp 1711653199
transform 1 0 1236 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3680
timestamp 1711653199
transform 1 0 1876 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3681
timestamp 1711653199
transform 1 0 1796 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3682
timestamp 1711653199
transform 1 0 2060 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3683
timestamp 1711653199
transform 1 0 1836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3684
timestamp 1711653199
transform 1 0 2652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3685
timestamp 1711653199
transform 1 0 2636 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1711653199
transform 1 0 2012 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3687
timestamp 1711653199
transform 1 0 2036 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3688
timestamp 1711653199
transform 1 0 2028 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3689
timestamp 1711653199
transform 1 0 2164 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3690
timestamp 1711653199
transform 1 0 2140 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1711653199
transform 1 0 1980 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3692
timestamp 1711653199
transform 1 0 1900 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_3693
timestamp 1711653199
transform 1 0 2180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3694
timestamp 1711653199
transform 1 0 2172 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3695
timestamp 1711653199
transform 1 0 1844 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3696
timestamp 1711653199
transform 1 0 1684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_3697
timestamp 1711653199
transform 1 0 1876 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3698
timestamp 1711653199
transform 1 0 1876 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3699
timestamp 1711653199
transform 1 0 1812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3700
timestamp 1711653199
transform 1 0 796 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3701
timestamp 1711653199
transform 1 0 748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3702
timestamp 1711653199
transform 1 0 748 0 1 1055
box -2 -2 2 2
use M2_M1  M2_M1_3703
timestamp 1711653199
transform 1 0 732 0 1 1055
box -2 -2 2 2
use M2_M1  M2_M1_3704
timestamp 1711653199
transform 1 0 700 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3705
timestamp 1711653199
transform 1 0 2276 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3706
timestamp 1711653199
transform 1 0 2244 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3707
timestamp 1711653199
transform 1 0 2244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3708
timestamp 1711653199
transform 1 0 1940 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3709
timestamp 1711653199
transform 1 0 1492 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3710
timestamp 1711653199
transform 1 0 740 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3711
timestamp 1711653199
transform 1 0 1644 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3712
timestamp 1711653199
transform 1 0 1548 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3713
timestamp 1711653199
transform 1 0 1852 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3714
timestamp 1711653199
transform 1 0 1692 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3715
timestamp 1711653199
transform 1 0 1716 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3716
timestamp 1711653199
transform 1 0 1492 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3717
timestamp 1711653199
transform 1 0 1924 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3718
timestamp 1711653199
transform 1 0 1788 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3719
timestamp 1711653199
transform 1 0 2148 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3720
timestamp 1711653199
transform 1 0 1980 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3721
timestamp 1711653199
transform 1 0 1900 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3722
timestamp 1711653199
transform 1 0 1924 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3723
timestamp 1711653199
transform 1 0 852 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3724
timestamp 1711653199
transform 1 0 3188 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3725
timestamp 1711653199
transform 1 0 2924 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3726
timestamp 1711653199
transform 1 0 2884 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3727
timestamp 1711653199
transform 1 0 2316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3728
timestamp 1711653199
transform 1 0 900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3729
timestamp 1711653199
transform 1 0 836 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3730
timestamp 1711653199
transform 1 0 916 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3731
timestamp 1711653199
transform 1 0 844 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3732
timestamp 1711653199
transform 1 0 860 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3733
timestamp 1711653199
transform 1 0 740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3734
timestamp 1711653199
transform 1 0 676 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3735
timestamp 1711653199
transform 1 0 1452 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3736
timestamp 1711653199
transform 1 0 852 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3737
timestamp 1711653199
transform 1 0 588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1711653199
transform 1 0 2484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3739
timestamp 1711653199
transform 1 0 2228 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_3740
timestamp 1711653199
transform 1 0 2172 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_3741
timestamp 1711653199
transform 1 0 2108 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_3742
timestamp 1711653199
transform 1 0 1468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3743
timestamp 1711653199
transform 1 0 1468 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3744
timestamp 1711653199
transform 1 0 1252 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3745
timestamp 1711653199
transform 1 0 1252 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_3746
timestamp 1711653199
transform 1 0 1004 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3747
timestamp 1711653199
transform 1 0 996 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_3748
timestamp 1711653199
transform 1 0 1516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3749
timestamp 1711653199
transform 1 0 1508 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3750
timestamp 1711653199
transform 1 0 1444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3751
timestamp 1711653199
transform 1 0 1428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3752
timestamp 1711653199
transform 1 0 652 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3753
timestamp 1711653199
transform 1 0 612 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_3754
timestamp 1711653199
transform 1 0 572 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3755
timestamp 1711653199
transform 1 0 1700 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3756
timestamp 1711653199
transform 1 0 1668 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3757
timestamp 1711653199
transform 1 0 1492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3758
timestamp 1711653199
transform 1 0 1524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3759
timestamp 1711653199
transform 1 0 1340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3760
timestamp 1711653199
transform 1 0 1324 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3761
timestamp 1711653199
transform 1 0 1924 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3762
timestamp 1711653199
transform 1 0 1892 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3763
timestamp 1711653199
transform 1 0 2556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3764
timestamp 1711653199
transform 1 0 1948 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3765
timestamp 1711653199
transform 1 0 2892 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3766
timestamp 1711653199
transform 1 0 2836 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3767
timestamp 1711653199
transform 1 0 2532 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3768
timestamp 1711653199
transform 1 0 2076 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3769
timestamp 1711653199
transform 1 0 2004 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3770
timestamp 1711653199
transform 1 0 1908 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3771
timestamp 1711653199
transform 1 0 1884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3772
timestamp 1711653199
transform 1 0 1828 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_3773
timestamp 1711653199
transform 1 0 1932 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3774
timestamp 1711653199
transform 1 0 1820 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3775
timestamp 1711653199
transform 1 0 2252 0 1 145
box -2 -2 2 2
use M2_M1  M2_M1_3776
timestamp 1711653199
transform 1 0 2236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3777
timestamp 1711653199
transform 1 0 2196 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3778
timestamp 1711653199
transform 1 0 2060 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1711653199
transform 1 0 1804 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3780
timestamp 1711653199
transform 1 0 1804 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3781
timestamp 1711653199
transform 1 0 252 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3782
timestamp 1711653199
transform 1 0 204 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3783
timestamp 1711653199
transform 1 0 1836 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3784
timestamp 1711653199
transform 1 0 1796 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3785
timestamp 1711653199
transform 1 0 1940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3786
timestamp 1711653199
transform 1 0 1924 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3787
timestamp 1711653199
transform 1 0 1892 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3788
timestamp 1711653199
transform 1 0 1892 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3789
timestamp 1711653199
transform 1 0 780 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3790
timestamp 1711653199
transform 1 0 684 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3791
timestamp 1711653199
transform 1 0 700 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_3792
timestamp 1711653199
transform 1 0 596 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3793
timestamp 1711653199
transform 1 0 548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3794
timestamp 1711653199
transform 1 0 548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3795
timestamp 1711653199
transform 1 0 500 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3796
timestamp 1711653199
transform 1 0 492 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3797
timestamp 1711653199
transform 1 0 492 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3798
timestamp 1711653199
transform 1 0 524 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3799
timestamp 1711653199
transform 1 0 196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3800
timestamp 1711653199
transform 1 0 204 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3801
timestamp 1711653199
transform 1 0 188 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3802
timestamp 1711653199
transform 1 0 188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3803
timestamp 1711653199
transform 1 0 236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3804
timestamp 1711653199
transform 1 0 196 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3805
timestamp 1711653199
transform 1 0 164 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3806
timestamp 1711653199
transform 1 0 1668 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3807
timestamp 1711653199
transform 1 0 524 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3808
timestamp 1711653199
transform 1 0 2972 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3809
timestamp 1711653199
transform 1 0 1660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3810
timestamp 1711653199
transform 1 0 1676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3811
timestamp 1711653199
transform 1 0 1348 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3812
timestamp 1711653199
transform 1 0 1324 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3813
timestamp 1711653199
transform 1 0 2916 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3814
timestamp 1711653199
transform 1 0 2916 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3815
timestamp 1711653199
transform 1 0 3124 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3816
timestamp 1711653199
transform 1 0 3020 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3817
timestamp 1711653199
transform 1 0 3236 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3818
timestamp 1711653199
transform 1 0 3228 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3819
timestamp 1711653199
transform 1 0 3116 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3820
timestamp 1711653199
transform 1 0 3220 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3821
timestamp 1711653199
transform 1 0 3156 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3822
timestamp 1711653199
transform 1 0 3156 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1711653199
transform 1 0 412 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3824
timestamp 1711653199
transform 1 0 300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3825
timestamp 1711653199
transform 1 0 852 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3826
timestamp 1711653199
transform 1 0 764 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_3827
timestamp 1711653199
transform 1 0 820 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3828
timestamp 1711653199
transform 1 0 812 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3829
timestamp 1711653199
transform 1 0 764 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3830
timestamp 1711653199
transform 1 0 764 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3831
timestamp 1711653199
transform 1 0 1284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3832
timestamp 1711653199
transform 1 0 844 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3833
timestamp 1711653199
transform 1 0 1468 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3834
timestamp 1711653199
transform 1 0 1452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3835
timestamp 1711653199
transform 1 0 1252 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3836
timestamp 1711653199
transform 1 0 548 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3837
timestamp 1711653199
transform 1 0 252 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_3838
timestamp 1711653199
transform 1 0 236 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3839
timestamp 1711653199
transform 1 0 1580 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_3840
timestamp 1711653199
transform 1 0 1580 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3841
timestamp 1711653199
transform 1 0 1276 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3842
timestamp 1711653199
transform 1 0 1300 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3843
timestamp 1711653199
transform 1 0 1252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3844
timestamp 1711653199
transform 1 0 796 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1711653199
transform 1 0 756 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3846
timestamp 1711653199
transform 1 0 900 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3847
timestamp 1711653199
transform 1 0 860 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3848
timestamp 1711653199
transform 1 0 860 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3849
timestamp 1711653199
transform 1 0 380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3850
timestamp 1711653199
transform 1 0 268 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3851
timestamp 1711653199
transform 1 0 1100 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3852
timestamp 1711653199
transform 1 0 948 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3853
timestamp 1711653199
transform 1 0 1420 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3854
timestamp 1711653199
transform 1 0 1420 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3855
timestamp 1711653199
transform 1 0 1476 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3856
timestamp 1711653199
transform 1 0 1468 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3857
timestamp 1711653199
transform 1 0 1932 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3858
timestamp 1711653199
transform 1 0 1500 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3859
timestamp 1711653199
transform 1 0 1532 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3860
timestamp 1711653199
transform 1 0 1532 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3861
timestamp 1711653199
transform 1 0 1572 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3862
timestamp 1711653199
transform 1 0 1524 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3863
timestamp 1711653199
transform 1 0 1540 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3864
timestamp 1711653199
transform 1 0 852 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3865
timestamp 1711653199
transform 1 0 820 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3866
timestamp 1711653199
transform 1 0 732 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3867
timestamp 1711653199
transform 1 0 676 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3868
timestamp 1711653199
transform 1 0 2364 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3869
timestamp 1711653199
transform 1 0 2068 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3870
timestamp 1711653199
transform 1 0 1740 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3871
timestamp 1711653199
transform 1 0 884 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3872
timestamp 1711653199
transform 1 0 812 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3873
timestamp 1711653199
transform 1 0 660 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_3874
timestamp 1711653199
transform 1 0 468 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_3875
timestamp 1711653199
transform 1 0 444 0 1 1245
box -2 -2 2 2
use M2_M1  M2_M1_3876
timestamp 1711653199
transform 1 0 388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_3877
timestamp 1711653199
transform 1 0 340 0 1 845
box -2 -2 2 2
use M2_M1  M2_M1_3878
timestamp 1711653199
transform 1 0 332 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_3879
timestamp 1711653199
transform 1 0 300 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_3880
timestamp 1711653199
transform 1 0 884 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3881
timestamp 1711653199
transform 1 0 860 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3882
timestamp 1711653199
transform 1 0 876 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3883
timestamp 1711653199
transform 1 0 860 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3884
timestamp 1711653199
transform 1 0 860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3885
timestamp 1711653199
transform 1 0 852 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3886
timestamp 1711653199
transform 1 0 892 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3887
timestamp 1711653199
transform 1 0 844 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3888
timestamp 1711653199
transform 1 0 844 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3889
timestamp 1711653199
transform 1 0 1500 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3890
timestamp 1711653199
transform 1 0 1236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3891
timestamp 1711653199
transform 1 0 1572 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3892
timestamp 1711653199
transform 1 0 1412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3893
timestamp 1711653199
transform 1 0 1404 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3894
timestamp 1711653199
transform 1 0 692 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3895
timestamp 1711653199
transform 1 0 692 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3896
timestamp 1711653199
transform 1 0 1684 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3897
timestamp 1711653199
transform 1 0 1572 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3898
timestamp 1711653199
transform 1 0 1468 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3899
timestamp 1711653199
transform 1 0 2036 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3900
timestamp 1711653199
transform 1 0 1956 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_3901
timestamp 1711653199
transform 1 0 2108 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3902
timestamp 1711653199
transform 1 0 1996 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_3903
timestamp 1711653199
transform 1 0 2068 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3904
timestamp 1711653199
transform 1 0 2028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_3905
timestamp 1711653199
transform 1 0 1940 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_3906
timestamp 1711653199
transform 1 0 2596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3907
timestamp 1711653199
transform 1 0 2564 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3908
timestamp 1711653199
transform 1 0 2604 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3909
timestamp 1711653199
transform 1 0 2572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3910
timestamp 1711653199
transform 1 0 2564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_3911
timestamp 1711653199
transform 1 0 2532 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3912
timestamp 1711653199
transform 1 0 2588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3913
timestamp 1711653199
transform 1 0 2444 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3914
timestamp 1711653199
transform 1 0 2476 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_3915
timestamp 1711653199
transform 1 0 2380 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_3916
timestamp 1711653199
transform 1 0 2380 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_3917
timestamp 1711653199
transform 1 0 2156 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_3918
timestamp 1711653199
transform 1 0 2516 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3919
timestamp 1711653199
transform 1 0 2460 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3920
timestamp 1711653199
transform 1 0 2356 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3921
timestamp 1711653199
transform 1 0 2356 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_3922
timestamp 1711653199
transform 1 0 2596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_3923
timestamp 1711653199
transform 1 0 2580 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_3924
timestamp 1711653199
transform 1 0 2508 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_3925
timestamp 1711653199
transform 1 0 2404 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_3926
timestamp 1711653199
transform 1 0 2060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3927
timestamp 1711653199
transform 1 0 1988 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3928
timestamp 1711653199
transform 1 0 1988 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3929
timestamp 1711653199
transform 1 0 2044 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3930
timestamp 1711653199
transform 1 0 2044 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3931
timestamp 1711653199
transform 1 0 2180 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3932
timestamp 1711653199
transform 1 0 2164 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3933
timestamp 1711653199
transform 1 0 2036 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3934
timestamp 1711653199
transform 1 0 2060 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_3935
timestamp 1711653199
transform 1 0 1804 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3936
timestamp 1711653199
transform 1 0 1804 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_3937
timestamp 1711653199
transform 1 0 1412 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3938
timestamp 1711653199
transform 1 0 1412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3939
timestamp 1711653199
transform 1 0 1604 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3940
timestamp 1711653199
transform 1 0 1460 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_3941
timestamp 1711653199
transform 1 0 1476 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3942
timestamp 1711653199
transform 1 0 124 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3943
timestamp 1711653199
transform 1 0 124 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3944
timestamp 1711653199
transform 1 0 108 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3945
timestamp 1711653199
transform 1 0 308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3946
timestamp 1711653199
transform 1 0 164 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3947
timestamp 1711653199
transform 1 0 100 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3948
timestamp 1711653199
transform 1 0 148 0 1 385
box -2 -2 2 2
use M2_M1  M2_M1_3949
timestamp 1711653199
transform 1 0 148 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3950
timestamp 1711653199
transform 1 0 132 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3951
timestamp 1711653199
transform 1 0 108 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3952
timestamp 1711653199
transform 1 0 100 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3953
timestamp 1711653199
transform 1 0 92 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3954
timestamp 1711653199
transform 1 0 92 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3955
timestamp 1711653199
transform 1 0 2852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3956
timestamp 1711653199
transform 1 0 1644 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_3957
timestamp 1711653199
transform 1 0 2860 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3958
timestamp 1711653199
transform 1 0 2852 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3959
timestamp 1711653199
transform 1 0 2844 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3960
timestamp 1711653199
transform 1 0 3068 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3961
timestamp 1711653199
transform 1 0 2908 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3962
timestamp 1711653199
transform 1 0 3084 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_3963
timestamp 1711653199
transform 1 0 3084 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3964
timestamp 1711653199
transform 1 0 3044 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3965
timestamp 1711653199
transform 1 0 3212 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3966
timestamp 1711653199
transform 1 0 3100 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_3967
timestamp 1711653199
transform 1 0 3276 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3968
timestamp 1711653199
transform 1 0 3268 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3969
timestamp 1711653199
transform 1 0 3204 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3970
timestamp 1711653199
transform 1 0 3204 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_3971
timestamp 1711653199
transform 1 0 3276 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_3972
timestamp 1711653199
transform 1 0 3260 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_3973
timestamp 1711653199
transform 1 0 3252 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_3974
timestamp 1711653199
transform 1 0 1516 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3975
timestamp 1711653199
transform 1 0 1500 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_3976
timestamp 1711653199
transform 1 0 1364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3977
timestamp 1711653199
transform 1 0 1340 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_3978
timestamp 1711653199
transform 1 0 1372 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3979
timestamp 1711653199
transform 1 0 1372 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_3980
timestamp 1711653199
transform 1 0 1444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3981
timestamp 1711653199
transform 1 0 1444 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_3982
timestamp 1711653199
transform 1 0 1380 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3983
timestamp 1711653199
transform 1 0 1228 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3984
timestamp 1711653199
transform 1 0 1188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3985
timestamp 1711653199
transform 1 0 1452 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3986
timestamp 1711653199
transform 1 0 1452 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3987
timestamp 1711653199
transform 1 0 1404 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3988
timestamp 1711653199
transform 1 0 1004 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3989
timestamp 1711653199
transform 1 0 980 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3990
timestamp 1711653199
transform 1 0 1740 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3991
timestamp 1711653199
transform 1 0 1532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_3992
timestamp 1711653199
transform 1 0 1500 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_3993
timestamp 1711653199
transform 1 0 1500 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_3994
timestamp 1711653199
transform 1 0 1324 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3995
timestamp 1711653199
transform 1 0 1116 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_3996
timestamp 1711653199
transform 1 0 932 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_3997
timestamp 1711653199
transform 1 0 1372 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_3998
timestamp 1711653199
transform 1 0 492 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_3999
timestamp 1711653199
transform 1 0 444 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4000
timestamp 1711653199
transform 1 0 380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4001
timestamp 1711653199
transform 1 0 348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4002
timestamp 1711653199
transform 1 0 500 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4003
timestamp 1711653199
transform 1 0 220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4004
timestamp 1711653199
transform 1 0 212 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4005
timestamp 1711653199
transform 1 0 2196 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4006
timestamp 1711653199
transform 1 0 2180 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4007
timestamp 1711653199
transform 1 0 2396 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4008
timestamp 1711653199
transform 1 0 2164 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4009
timestamp 1711653199
transform 1 0 2156 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4010
timestamp 1711653199
transform 1 0 2156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4011
timestamp 1711653199
transform 1 0 2156 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4012
timestamp 1711653199
transform 1 0 2100 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4013
timestamp 1711653199
transform 1 0 2156 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4014
timestamp 1711653199
transform 1 0 2012 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4015
timestamp 1711653199
transform 1 0 1996 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4016
timestamp 1711653199
transform 1 0 1996 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4017
timestamp 1711653199
transform 1 0 2428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4018
timestamp 1711653199
transform 1 0 2412 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4019
timestamp 1711653199
transform 1 0 2748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4020
timestamp 1711653199
transform 1 0 2540 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4021
timestamp 1711653199
transform 1 0 2484 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4022
timestamp 1711653199
transform 1 0 2412 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4023
timestamp 1711653199
transform 1 0 2388 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4024
timestamp 1711653199
transform 1 0 2388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4025
timestamp 1711653199
transform 1 0 2108 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4026
timestamp 1711653199
transform 1 0 2036 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4027
timestamp 1711653199
transform 1 0 2004 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4028
timestamp 1711653199
transform 1 0 2356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4029
timestamp 1711653199
transform 1 0 2332 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4030
timestamp 1711653199
transform 1 0 2140 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4031
timestamp 1711653199
transform 1 0 2132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4032
timestamp 1711653199
transform 1 0 2060 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4033
timestamp 1711653199
transform 1 0 2004 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4034
timestamp 1711653199
transform 1 0 1996 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4035
timestamp 1711653199
transform 1 0 1980 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4036
timestamp 1711653199
transform 1 0 1980 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4037
timestamp 1711653199
transform 1 0 1972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4038
timestamp 1711653199
transform 1 0 1748 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_4039
timestamp 1711653199
transform 1 0 2140 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4040
timestamp 1711653199
transform 1 0 2084 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4041
timestamp 1711653199
transform 1 0 2164 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4042
timestamp 1711653199
transform 1 0 2108 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4043
timestamp 1711653199
transform 1 0 2252 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4044
timestamp 1711653199
transform 1 0 2092 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4045
timestamp 1711653199
transform 1 0 2484 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4046
timestamp 1711653199
transform 1 0 2228 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4047
timestamp 1711653199
transform 1 0 2252 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4048
timestamp 1711653199
transform 1 0 2236 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4049
timestamp 1711653199
transform 1 0 2268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4050
timestamp 1711653199
transform 1 0 2252 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4051
timestamp 1711653199
transform 1 0 2364 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4052
timestamp 1711653199
transform 1 0 2324 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4053
timestamp 1711653199
transform 1 0 2196 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4054
timestamp 1711653199
transform 1 0 2092 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4055
timestamp 1711653199
transform 1 0 2500 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4056
timestamp 1711653199
transform 1 0 2476 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4057
timestamp 1711653199
transform 1 0 2444 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4058
timestamp 1711653199
transform 1 0 2420 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4059
timestamp 1711653199
transform 1 0 2396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4060
timestamp 1711653199
transform 1 0 2156 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4061
timestamp 1711653199
transform 1 0 1900 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4062
timestamp 1711653199
transform 1 0 2052 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4063
timestamp 1711653199
transform 1 0 2020 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4064
timestamp 1711653199
transform 1 0 1636 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4065
timestamp 1711653199
transform 1 0 1636 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_4066
timestamp 1711653199
transform 1 0 2284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4067
timestamp 1711653199
transform 1 0 2052 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4068
timestamp 1711653199
transform 1 0 2508 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4069
timestamp 1711653199
transform 1 0 2260 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4070
timestamp 1711653199
transform 1 0 2292 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4071
timestamp 1711653199
transform 1 0 2260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4072
timestamp 1711653199
transform 1 0 2324 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_4073
timestamp 1711653199
transform 1 0 2324 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4074
timestamp 1711653199
transform 1 0 2388 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4075
timestamp 1711653199
transform 1 0 2356 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4076
timestamp 1711653199
transform 1 0 2228 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4077
timestamp 1711653199
transform 1 0 2108 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4078
timestamp 1711653199
transform 1 0 2588 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4079
timestamp 1711653199
transform 1 0 2540 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4080
timestamp 1711653199
transform 1 0 2596 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4081
timestamp 1711653199
transform 1 0 2516 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4082
timestamp 1711653199
transform 1 0 2500 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4083
timestamp 1711653199
transform 1 0 2156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4084
timestamp 1711653199
transform 1 0 2156 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4085
timestamp 1711653199
transform 1 0 3172 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4086
timestamp 1711653199
transform 1 0 3156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4087
timestamp 1711653199
transform 1 0 2836 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4088
timestamp 1711653199
transform 1 0 2780 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_4089
timestamp 1711653199
transform 1 0 2908 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4090
timestamp 1711653199
transform 1 0 2868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4091
timestamp 1711653199
transform 1 0 2836 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4092
timestamp 1711653199
transform 1 0 2716 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4093
timestamp 1711653199
transform 1 0 2652 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4094
timestamp 1711653199
transform 1 0 2060 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4095
timestamp 1711653199
transform 1 0 1932 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4096
timestamp 1711653199
transform 1 0 2252 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4097
timestamp 1711653199
transform 1 0 2028 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4098
timestamp 1711653199
transform 1 0 2012 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4099
timestamp 1711653199
transform 1 0 1980 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4100
timestamp 1711653199
transform 1 0 1940 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4101
timestamp 1711653199
transform 1 0 1916 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4102
timestamp 1711653199
transform 1 0 2012 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4103
timestamp 1711653199
transform 1 0 1964 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4104
timestamp 1711653199
transform 1 0 1964 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4105
timestamp 1711653199
transform 1 0 1948 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4106
timestamp 1711653199
transform 1 0 1932 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4107
timestamp 1711653199
transform 1 0 2116 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4108
timestamp 1711653199
transform 1 0 2076 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4109
timestamp 1711653199
transform 1 0 2172 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4110
timestamp 1711653199
transform 1 0 2116 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4111
timestamp 1711653199
transform 1 0 2356 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4112
timestamp 1711653199
transform 1 0 2220 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4113
timestamp 1711653199
transform 1 0 2132 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4114
timestamp 1711653199
transform 1 0 2132 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4115
timestamp 1711653199
transform 1 0 2116 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4116
timestamp 1711653199
transform 1 0 2100 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4117
timestamp 1711653199
transform 1 0 2420 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4118
timestamp 1711653199
transform 1 0 2380 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4119
timestamp 1711653199
transform 1 0 2340 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4120
timestamp 1711653199
transform 1 0 2148 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4121
timestamp 1711653199
transform 1 0 2132 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4122
timestamp 1711653199
transform 1 0 2100 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4123
timestamp 1711653199
transform 1 0 2460 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4124
timestamp 1711653199
transform 1 0 2412 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4125
timestamp 1711653199
transform 1 0 2236 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4126
timestamp 1711653199
transform 1 0 2092 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4127
timestamp 1711653199
transform 1 0 1964 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4128
timestamp 1711653199
transform 1 0 1636 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4129
timestamp 1711653199
transform 1 0 1612 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4130
timestamp 1711653199
transform 1 0 1524 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4131
timestamp 1711653199
transform 1 0 2300 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4132
timestamp 1711653199
transform 1 0 2276 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_4133
timestamp 1711653199
transform 1 0 2124 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4134
timestamp 1711653199
transform 1 0 2060 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4135
timestamp 1711653199
transform 1 0 1772 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4136
timestamp 1711653199
transform 1 0 1668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4137
timestamp 1711653199
transform 1 0 1652 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4138
timestamp 1711653199
transform 1 0 1620 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_4139
timestamp 1711653199
transform 1 0 2332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4140
timestamp 1711653199
transform 1 0 2284 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4141
timestamp 1711653199
transform 1 0 2404 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4142
timestamp 1711653199
transform 1 0 2308 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4143
timestamp 1711653199
transform 1 0 2356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4144
timestamp 1711653199
transform 1 0 2188 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4145
timestamp 1711653199
transform 1 0 2148 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4146
timestamp 1711653199
transform 1 0 2196 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4147
timestamp 1711653199
transform 1 0 2116 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4148
timestamp 1711653199
transform 1 0 2108 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4149
timestamp 1711653199
transform 1 0 2020 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4150
timestamp 1711653199
transform 1 0 1964 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4151
timestamp 1711653199
transform 1 0 1868 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4152
timestamp 1711653199
transform 1 0 1820 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4153
timestamp 1711653199
transform 1 0 1580 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4154
timestamp 1711653199
transform 1 0 1516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4155
timestamp 1711653199
transform 1 0 1444 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4156
timestamp 1711653199
transform 1 0 1068 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_4157
timestamp 1711653199
transform 1 0 1044 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4158
timestamp 1711653199
transform 1 0 1996 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4159
timestamp 1711653199
transform 1 0 1596 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4160
timestamp 1711653199
transform 1 0 1596 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4161
timestamp 1711653199
transform 1 0 1100 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4162
timestamp 1711653199
transform 1 0 1052 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4163
timestamp 1711653199
transform 1 0 732 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4164
timestamp 1711653199
transform 1 0 2108 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4165
timestamp 1711653199
transform 1 0 2044 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4166
timestamp 1711653199
transform 1 0 2020 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4167
timestamp 1711653199
transform 1 0 1956 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4168
timestamp 1711653199
transform 1 0 1900 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4169
timestamp 1711653199
transform 1 0 2204 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4170
timestamp 1711653199
transform 1 0 2204 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4171
timestamp 1711653199
transform 1 0 1796 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4172
timestamp 1711653199
transform 1 0 1684 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4173
timestamp 1711653199
transform 1 0 2020 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4174
timestamp 1711653199
transform 1 0 1772 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4175
timestamp 1711653199
transform 1 0 1900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4176
timestamp 1711653199
transform 1 0 1780 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4177
timestamp 1711653199
transform 1 0 1884 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4178
timestamp 1711653199
transform 1 0 1868 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4179
timestamp 1711653199
transform 1 0 1980 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4180
timestamp 1711653199
transform 1 0 1924 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4181
timestamp 1711653199
transform 1 0 2044 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4182
timestamp 1711653199
transform 1 0 2044 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4183
timestamp 1711653199
transform 1 0 1908 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4184
timestamp 1711653199
transform 1 0 2348 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4185
timestamp 1711653199
transform 1 0 2156 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4186
timestamp 1711653199
transform 1 0 2068 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4187
timestamp 1711653199
transform 1 0 1996 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4188
timestamp 1711653199
transform 1 0 1812 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4189
timestamp 1711653199
transform 1 0 1308 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4190
timestamp 1711653199
transform 1 0 564 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4191
timestamp 1711653199
transform 1 0 308 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4192
timestamp 1711653199
transform 1 0 268 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4193
timestamp 1711653199
transform 1 0 252 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4194
timestamp 1711653199
transform 1 0 2132 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4195
timestamp 1711653199
transform 1 0 2132 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4196
timestamp 1711653199
transform 1 0 2124 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4197
timestamp 1711653199
transform 1 0 1892 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4198
timestamp 1711653199
transform 1 0 1788 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4199
timestamp 1711653199
transform 1 0 1740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4200
timestamp 1711653199
transform 1 0 1740 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4201
timestamp 1711653199
transform 1 0 1740 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4202
timestamp 1711653199
transform 1 0 1724 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4203
timestamp 1711653199
transform 1 0 932 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4204
timestamp 1711653199
transform 1 0 932 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_4205
timestamp 1711653199
transform 1 0 908 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_4206
timestamp 1711653199
transform 1 0 684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4207
timestamp 1711653199
transform 1 0 1788 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4208
timestamp 1711653199
transform 1 0 1764 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4209
timestamp 1711653199
transform 1 0 2372 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4210
timestamp 1711653199
transform 1 0 2332 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4211
timestamp 1711653199
transform 1 0 2220 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4212
timestamp 1711653199
transform 1 0 1940 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_4213
timestamp 1711653199
transform 1 0 1868 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4214
timestamp 1711653199
transform 1 0 884 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4215
timestamp 1711653199
transform 1 0 884 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4216
timestamp 1711653199
transform 1 0 2164 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4217
timestamp 1711653199
transform 1 0 1996 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4218
timestamp 1711653199
transform 1 0 2068 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4219
timestamp 1711653199
transform 1 0 2004 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4220
timestamp 1711653199
transform 1 0 2756 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4221
timestamp 1711653199
transform 1 0 2692 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4222
timestamp 1711653199
transform 1 0 2692 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4223
timestamp 1711653199
transform 1 0 2332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4224
timestamp 1711653199
transform 1 0 2180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4225
timestamp 1711653199
transform 1 0 2076 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4226
timestamp 1711653199
transform 1 0 1948 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4227
timestamp 1711653199
transform 1 0 1788 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4228
timestamp 1711653199
transform 1 0 1748 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4229
timestamp 1711653199
transform 1 0 1196 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4230
timestamp 1711653199
transform 1 0 1036 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4231
timestamp 1711653199
transform 1 0 1036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4232
timestamp 1711653199
transform 1 0 1004 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4233
timestamp 1711653199
transform 1 0 708 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4234
timestamp 1711653199
transform 1 0 580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4235
timestamp 1711653199
transform 1 0 564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4236
timestamp 1711653199
transform 1 0 500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4237
timestamp 1711653199
transform 1 0 2036 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4238
timestamp 1711653199
transform 1 0 2036 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4239
timestamp 1711653199
transform 1 0 3012 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4240
timestamp 1711653199
transform 1 0 2868 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4241
timestamp 1711653199
transform 1 0 2828 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4242
timestamp 1711653199
transform 1 0 2140 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4243
timestamp 1711653199
transform 1 0 2140 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4244
timestamp 1711653199
transform 1 0 2028 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_4245
timestamp 1711653199
transform 1 0 1300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4246
timestamp 1711653199
transform 1 0 1260 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4247
timestamp 1711653199
transform 1 0 964 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4248
timestamp 1711653199
transform 1 0 844 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4249
timestamp 1711653199
transform 1 0 780 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4250
timestamp 1711653199
transform 1 0 732 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4251
timestamp 1711653199
transform 1 0 2156 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4252
timestamp 1711653199
transform 1 0 2132 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4253
timestamp 1711653199
transform 1 0 2300 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4254
timestamp 1711653199
transform 1 0 1812 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4255
timestamp 1711653199
transform 1 0 1764 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4256
timestamp 1711653199
transform 1 0 908 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4257
timestamp 1711653199
transform 1 0 892 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4258
timestamp 1711653199
transform 1 0 2836 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4259
timestamp 1711653199
transform 1 0 2596 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4260
timestamp 1711653199
transform 1 0 2396 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4261
timestamp 1711653199
transform 1 0 2268 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_4262
timestamp 1711653199
transform 1 0 2244 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4263
timestamp 1711653199
transform 1 0 1844 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4264
timestamp 1711653199
transform 1 0 1796 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_4265
timestamp 1711653199
transform 1 0 1252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4266
timestamp 1711653199
transform 1 0 1004 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4267
timestamp 1711653199
transform 1 0 1884 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4268
timestamp 1711653199
transform 1 0 1812 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4269
timestamp 1711653199
transform 1 0 1580 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4270
timestamp 1711653199
transform 1 0 1524 0 1 1985
box -2 -2 2 2
use M2_M1  M2_M1_4271
timestamp 1711653199
transform 1 0 1484 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4272
timestamp 1711653199
transform 1 0 1484 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_4273
timestamp 1711653199
transform 1 0 1604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4274
timestamp 1711653199
transform 1 0 1540 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4275
timestamp 1711653199
transform 1 0 1708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4276
timestamp 1711653199
transform 1 0 1548 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4277
timestamp 1711653199
transform 1 0 1724 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4278
timestamp 1711653199
transform 1 0 1676 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4279
timestamp 1711653199
transform 1 0 1900 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4280
timestamp 1711653199
transform 1 0 1748 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4281
timestamp 1711653199
transform 1 0 2228 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4282
timestamp 1711653199
transform 1 0 1964 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4283
timestamp 1711653199
transform 1 0 1892 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4284
timestamp 1711653199
transform 1 0 1892 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4285
timestamp 1711653199
transform 1 0 1604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4286
timestamp 1711653199
transform 1 0 1300 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4287
timestamp 1711653199
transform 1 0 236 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4288
timestamp 1711653199
transform 1 0 108 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4289
timestamp 1711653199
transform 1 0 108 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4290
timestamp 1711653199
transform 1 0 1908 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4291
timestamp 1711653199
transform 1 0 1900 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4292
timestamp 1711653199
transform 1 0 1716 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4293
timestamp 1711653199
transform 1 0 1708 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4294
timestamp 1711653199
transform 1 0 1684 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4295
timestamp 1711653199
transform 1 0 1628 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4296
timestamp 1711653199
transform 1 0 1716 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4297
timestamp 1711653199
transform 1 0 1684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4298
timestamp 1711653199
transform 1 0 1588 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4299
timestamp 1711653199
transform 1 0 1516 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4300
timestamp 1711653199
transform 1 0 1372 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4301
timestamp 1711653199
transform 1 0 1708 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4302
timestamp 1711653199
transform 1 0 1708 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4303
timestamp 1711653199
transform 1 0 1636 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4304
timestamp 1711653199
transform 1 0 1636 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4305
timestamp 1711653199
transform 1 0 1596 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4306
timestamp 1711653199
transform 1 0 1620 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4307
timestamp 1711653199
transform 1 0 1612 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_4308
timestamp 1711653199
transform 1 0 1660 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4309
timestamp 1711653199
transform 1 0 1548 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4310
timestamp 1711653199
transform 1 0 1156 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4311
timestamp 1711653199
transform 1 0 604 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4312
timestamp 1711653199
transform 1 0 2484 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4313
timestamp 1711653199
transform 1 0 2452 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4314
timestamp 1711653199
transform 1 0 2100 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4315
timestamp 1711653199
transform 1 0 2044 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4316
timestamp 1711653199
transform 1 0 1588 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_4317
timestamp 1711653199
transform 1 0 1108 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_4318
timestamp 1711653199
transform 1 0 1108 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_4319
timestamp 1711653199
transform 1 0 1108 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_4320
timestamp 1711653199
transform 1 0 1652 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4321
timestamp 1711653199
transform 1 0 1636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4322
timestamp 1711653199
transform 1 0 1964 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4323
timestamp 1711653199
transform 1 0 1780 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4324
timestamp 1711653199
transform 1 0 2028 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4325
timestamp 1711653199
transform 1 0 1988 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4326
timestamp 1711653199
transform 1 0 2436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4327
timestamp 1711653199
transform 1 0 1716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4328
timestamp 1711653199
transform 1 0 1572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4329
timestamp 1711653199
transform 1 0 1532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4330
timestamp 1711653199
transform 1 0 1276 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4331
timestamp 1711653199
transform 1 0 812 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4332
timestamp 1711653199
transform 1 0 2932 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4333
timestamp 1711653199
transform 1 0 2804 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4334
timestamp 1711653199
transform 1 0 2644 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4335
timestamp 1711653199
transform 1 0 2404 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4336
timestamp 1711653199
transform 1 0 1556 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4337
timestamp 1711653199
transform 1 0 1500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4338
timestamp 1711653199
transform 1 0 1732 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4339
timestamp 1711653199
transform 1 0 1692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4340
timestamp 1711653199
transform 1 0 1228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4341
timestamp 1711653199
transform 1 0 812 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4342
timestamp 1711653199
transform 1 0 1300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4343
timestamp 1711653199
transform 1 0 1260 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4344
timestamp 1711653199
transform 1 0 964 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4345
timestamp 1711653199
transform 1 0 772 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4346
timestamp 1711653199
transform 1 0 676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4347
timestamp 1711653199
transform 1 0 1572 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4348
timestamp 1711653199
transform 1 0 1324 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4349
timestamp 1711653199
transform 1 0 1564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4350
timestamp 1711653199
transform 1 0 1548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4351
timestamp 1711653199
transform 1 0 1612 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4352
timestamp 1711653199
transform 1 0 1548 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4353
timestamp 1711653199
transform 1 0 1636 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4354
timestamp 1711653199
transform 1 0 1636 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4355
timestamp 1711653199
transform 1 0 1756 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4356
timestamp 1711653199
transform 1 0 1740 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4357
timestamp 1711653199
transform 1 0 1684 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4358
timestamp 1711653199
transform 1 0 1684 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4359
timestamp 1711653199
transform 1 0 1852 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_4360
timestamp 1711653199
transform 1 0 1836 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4361
timestamp 1711653199
transform 1 0 1820 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4362
timestamp 1711653199
transform 1 0 1708 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4363
timestamp 1711653199
transform 1 0 1164 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4364
timestamp 1711653199
transform 1 0 404 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4365
timestamp 1711653199
transform 1 0 340 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4366
timestamp 1711653199
transform 1 0 316 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4367
timestamp 1711653199
transform 1 0 172 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4368
timestamp 1711653199
transform 1 0 1796 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_4369
timestamp 1711653199
transform 1 0 1788 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4370
timestamp 1711653199
transform 1 0 1668 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4371
timestamp 1711653199
transform 1 0 1636 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4372
timestamp 1711653199
transform 1 0 1556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4373
timestamp 1711653199
transform 1 0 1644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4374
timestamp 1711653199
transform 1 0 1644 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4375
timestamp 1711653199
transform 1 0 1588 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4376
timestamp 1711653199
transform 1 0 1452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4377
timestamp 1711653199
transform 1 0 1340 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4378
timestamp 1711653199
transform 1 0 1932 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4379
timestamp 1711653199
transform 1 0 1740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4380
timestamp 1711653199
transform 1 0 1708 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_4381
timestamp 1711653199
transform 1 0 1708 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4382
timestamp 1711653199
transform 1 0 1692 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_4383
timestamp 1711653199
transform 1 0 1692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4384
timestamp 1711653199
transform 1 0 1668 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4385
timestamp 1711653199
transform 1 0 1660 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_4386
timestamp 1711653199
transform 1 0 1628 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4387
timestamp 1711653199
transform 1 0 1516 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4388
timestamp 1711653199
transform 1 0 1244 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4389
timestamp 1711653199
transform 1 0 1052 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4390
timestamp 1711653199
transform 1 0 908 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4391
timestamp 1711653199
transform 1 0 1572 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4392
timestamp 1711653199
transform 1 0 1540 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4393
timestamp 1711653199
transform 1 0 1572 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4394
timestamp 1711653199
transform 1 0 1548 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4395
timestamp 1711653199
transform 1 0 1820 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4396
timestamp 1711653199
transform 1 0 1668 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4397
timestamp 1711653199
transform 1 0 1924 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4398
timestamp 1711653199
transform 1 0 1828 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4399
timestamp 1711653199
transform 1 0 2356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4400
timestamp 1711653199
transform 1 0 1484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4401
timestamp 1711653199
transform 1 0 1212 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4402
timestamp 1711653199
transform 1 0 1116 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4403
timestamp 1711653199
transform 1 0 876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4404
timestamp 1711653199
transform 1 0 2948 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4405
timestamp 1711653199
transform 1 0 2820 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4406
timestamp 1711653199
transform 1 0 2684 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4407
timestamp 1711653199
transform 1 0 2684 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_4408
timestamp 1711653199
transform 1 0 2420 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4409
timestamp 1711653199
transform 1 0 1532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4410
timestamp 1711653199
transform 1 0 1532 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4411
timestamp 1711653199
transform 1 0 1860 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4412
timestamp 1711653199
transform 1 0 1836 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4413
timestamp 1711653199
transform 1 0 1804 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4414
timestamp 1711653199
transform 1 0 1604 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4415
timestamp 1711653199
transform 1 0 1548 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4416
timestamp 1711653199
transform 1 0 1076 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4417
timestamp 1711653199
transform 1 0 1012 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4418
timestamp 1711653199
transform 1 0 1244 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4419
timestamp 1711653199
transform 1 0 1244 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4420
timestamp 1711653199
transform 1 0 972 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4421
timestamp 1711653199
transform 1 0 668 0 1 1985
box -2 -2 2 2
use M2_M1  M2_M1_4422
timestamp 1711653199
transform 1 0 652 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4423
timestamp 1711653199
transform 1 0 652 0 1 1985
box -2 -2 2 2
use M2_M1  M2_M1_4424
timestamp 1711653199
transform 1 0 300 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4425
timestamp 1711653199
transform 1 0 2028 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4426
timestamp 1711653199
transform 1 0 1148 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4427
timestamp 1711653199
transform 1 0 2028 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4428
timestamp 1711653199
transform 1 0 2004 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4429
timestamp 1711653199
transform 1 0 2028 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4430
timestamp 1711653199
transform 1 0 2012 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4431
timestamp 1711653199
transform 1 0 2044 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4432
timestamp 1711653199
transform 1 0 1940 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4433
timestamp 1711653199
transform 1 0 2140 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4434
timestamp 1711653199
transform 1 0 2116 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4435
timestamp 1711653199
transform 1 0 2116 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4436
timestamp 1711653199
transform 1 0 2084 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4437
timestamp 1711653199
transform 1 0 2044 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4438
timestamp 1711653199
transform 1 0 1948 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4439
timestamp 1711653199
transform 1 0 1916 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4440
timestamp 1711653199
transform 1 0 1596 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4441
timestamp 1711653199
transform 1 0 1156 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4442
timestamp 1711653199
transform 1 0 2116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4443
timestamp 1711653199
transform 1 0 2036 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4444
timestamp 1711653199
transform 1 0 1580 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_4445
timestamp 1711653199
transform 1 0 756 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4446
timestamp 1711653199
transform 1 0 2204 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4447
timestamp 1711653199
transform 1 0 2004 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_4448
timestamp 1711653199
transform 1 0 2020 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4449
timestamp 1711653199
transform 1 0 2012 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4450
timestamp 1711653199
transform 1 0 2196 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4451
timestamp 1711653199
transform 1 0 2188 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4452
timestamp 1711653199
transform 1 0 1852 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4453
timestamp 1711653199
transform 1 0 1844 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4454
timestamp 1711653199
transform 1 0 1860 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4455
timestamp 1711653199
transform 1 0 1860 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4456
timestamp 1711653199
transform 1 0 1644 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4457
timestamp 1711653199
transform 1 0 1044 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4458
timestamp 1711653199
transform 1 0 1044 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_4459
timestamp 1711653199
transform 1 0 1020 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_4460
timestamp 1711653199
transform 1 0 1012 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4461
timestamp 1711653199
transform 1 0 940 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4462
timestamp 1711653199
transform 1 0 1956 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4463
timestamp 1711653199
transform 1 0 1924 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4464
timestamp 1711653199
transform 1 0 1228 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4465
timestamp 1711653199
transform 1 0 1124 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4466
timestamp 1711653199
transform 1 0 876 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4467
timestamp 1711653199
transform 1 0 796 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4468
timestamp 1711653199
transform 1 0 788 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4469
timestamp 1711653199
transform 1 0 740 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4470
timestamp 1711653199
transform 1 0 1916 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4471
timestamp 1711653199
transform 1 0 1868 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4472
timestamp 1711653199
transform 1 0 2036 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4473
timestamp 1711653199
transform 1 0 1956 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4474
timestamp 1711653199
transform 1 0 1908 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4475
timestamp 1711653199
transform 1 0 1724 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4476
timestamp 1711653199
transform 1 0 484 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4477
timestamp 1711653199
transform 1 0 380 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4478
timestamp 1711653199
transform 1 0 532 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4479
timestamp 1711653199
transform 1 0 452 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4480
timestamp 1711653199
transform 1 0 604 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4481
timestamp 1711653199
transform 1 0 452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4482
timestamp 1711653199
transform 1 0 635 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4483
timestamp 1711653199
transform 1 0 612 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4484
timestamp 1711653199
transform 1 0 652 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4485
timestamp 1711653199
transform 1 0 652 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4486
timestamp 1711653199
transform 1 0 692 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4487
timestamp 1711653199
transform 1 0 668 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4488
timestamp 1711653199
transform 1 0 844 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4489
timestamp 1711653199
transform 1 0 668 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4490
timestamp 1711653199
transform 1 0 644 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4491
timestamp 1711653199
transform 1 0 628 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4492
timestamp 1711653199
transform 1 0 604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4493
timestamp 1711653199
transform 1 0 668 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4494
timestamp 1711653199
transform 1 0 628 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4495
timestamp 1711653199
transform 1 0 612 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4496
timestamp 1711653199
transform 1 0 612 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4497
timestamp 1711653199
transform 1 0 652 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_4498
timestamp 1711653199
transform 1 0 652 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4499
timestamp 1711653199
transform 1 0 1516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4500
timestamp 1711653199
transform 1 0 732 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4501
timestamp 1711653199
transform 1 0 628 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4502
timestamp 1711653199
transform 1 0 364 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4503
timestamp 1711653199
transform 1 0 620 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4504
timestamp 1711653199
transform 1 0 540 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_4505
timestamp 1711653199
transform 1 0 620 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4506
timestamp 1711653199
transform 1 0 596 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_4507
timestamp 1711653199
transform 1 0 2884 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4508
timestamp 1711653199
transform 1 0 2852 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4509
timestamp 1711653199
transform 1 0 2724 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4510
timestamp 1711653199
transform 1 0 2580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4511
timestamp 1711653199
transform 1 0 1964 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4512
timestamp 1711653199
transform 1 0 1852 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4513
timestamp 1711653199
transform 1 0 716 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4514
timestamp 1711653199
transform 1 0 708 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_4515
timestamp 1711653199
transform 1 0 684 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_4516
timestamp 1711653199
transform 1 0 628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4517
timestamp 1711653199
transform 1 0 692 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4518
timestamp 1711653199
transform 1 0 676 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4519
timestamp 1711653199
transform 1 0 700 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4520
timestamp 1711653199
transform 1 0 636 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4521
timestamp 1711653199
transform 1 0 564 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_4522
timestamp 1711653199
transform 1 0 556 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4523
timestamp 1711653199
transform 1 0 988 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4524
timestamp 1711653199
transform 1 0 708 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_4525
timestamp 1711653199
transform 1 0 2324 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4526
timestamp 1711653199
transform 1 0 2252 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4527
timestamp 1711653199
transform 1 0 2212 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4528
timestamp 1711653199
transform 1 0 1996 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_4529
timestamp 1711653199
transform 1 0 1900 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4530
timestamp 1711653199
transform 1 0 1596 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4531
timestamp 1711653199
transform 1 0 1588 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4532
timestamp 1711653199
transform 1 0 260 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4533
timestamp 1711653199
transform 1 0 124 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4534
timestamp 1711653199
transform 1 0 172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4535
timestamp 1711653199
transform 1 0 76 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_4536
timestamp 1711653199
transform 1 0 148 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4537
timestamp 1711653199
transform 1 0 108 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4538
timestamp 1711653199
transform 1 0 228 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4539
timestamp 1711653199
transform 1 0 124 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4540
timestamp 1711653199
transform 1 0 228 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4541
timestamp 1711653199
transform 1 0 180 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4542
timestamp 1711653199
transform 1 0 244 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4543
timestamp 1711653199
transform 1 0 244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4544
timestamp 1711653199
transform 1 0 348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4545
timestamp 1711653199
transform 1 0 316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4546
timestamp 1711653199
transform 1 0 228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4547
timestamp 1711653199
transform 1 0 172 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4548
timestamp 1711653199
transform 1 0 276 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4549
timestamp 1711653199
transform 1 0 244 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4550
timestamp 1711653199
transform 1 0 564 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4551
timestamp 1711653199
transform 1 0 548 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4552
timestamp 1711653199
transform 1 0 428 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4553
timestamp 1711653199
transform 1 0 412 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4554
timestamp 1711653199
transform 1 0 252 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_4555
timestamp 1711653199
transform 1 0 228 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4556
timestamp 1711653199
transform 1 0 196 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4557
timestamp 1711653199
transform 1 0 188 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4558
timestamp 1711653199
transform 1 0 188 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4559
timestamp 1711653199
transform 1 0 172 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4560
timestamp 1711653199
transform 1 0 220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4561
timestamp 1711653199
transform 1 0 204 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4562
timestamp 1711653199
transform 1 0 220 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4563
timestamp 1711653199
transform 1 0 204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4564
timestamp 1711653199
transform 1 0 188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4565
timestamp 1711653199
transform 1 0 188 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_4566
timestamp 1711653199
transform 1 0 244 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4567
timestamp 1711653199
transform 1 0 132 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4568
timestamp 1711653199
transform 1 0 212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4569
timestamp 1711653199
transform 1 0 188 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4570
timestamp 1711653199
transform 1 0 356 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4571
timestamp 1711653199
transform 1 0 340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4572
timestamp 1711653199
transform 1 0 332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4573
timestamp 1711653199
transform 1 0 468 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4574
timestamp 1711653199
transform 1 0 316 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4575
timestamp 1711653199
transform 1 0 348 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4576
timestamp 1711653199
transform 1 0 260 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4577
timestamp 1711653199
transform 1 0 284 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4578
timestamp 1711653199
transform 1 0 220 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4579
timestamp 1711653199
transform 1 0 860 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4580
timestamp 1711653199
transform 1 0 564 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4581
timestamp 1711653199
transform 1 0 532 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4582
timestamp 1711653199
transform 1 0 692 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4583
timestamp 1711653199
transform 1 0 460 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4584
timestamp 1711653199
transform 1 0 228 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4585
timestamp 1711653199
transform 1 0 108 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4586
timestamp 1711653199
transform 1 0 68 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4587
timestamp 1711653199
transform 1 0 68 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4588
timestamp 1711653199
transform 1 0 108 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4589
timestamp 1711653199
transform 1 0 92 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4590
timestamp 1711653199
transform 1 0 180 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4591
timestamp 1711653199
transform 1 0 116 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4592
timestamp 1711653199
transform 1 0 156 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4593
timestamp 1711653199
transform 1 0 148 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4594
timestamp 1711653199
transform 1 0 108 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4595
timestamp 1711653199
transform 1 0 92 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4596
timestamp 1711653199
transform 1 0 132 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4597
timestamp 1711653199
transform 1 0 108 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4598
timestamp 1711653199
transform 1 0 92 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4599
timestamp 1711653199
transform 1 0 92 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4600
timestamp 1711653199
transform 1 0 188 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4601
timestamp 1711653199
transform 1 0 116 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4602
timestamp 1711653199
transform 1 0 148 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4603
timestamp 1711653199
transform 1 0 116 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4604
timestamp 1711653199
transform 1 0 132 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4605
timestamp 1711653199
transform 1 0 132 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4606
timestamp 1711653199
transform 1 0 308 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4607
timestamp 1711653199
transform 1 0 276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4608
timestamp 1711653199
transform 1 0 220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4609
timestamp 1711653199
transform 1 0 116 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4610
timestamp 1711653199
transform 1 0 116 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4611
timestamp 1711653199
transform 1 0 108 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4612
timestamp 1711653199
transform 1 0 68 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4613
timestamp 1711653199
transform 1 0 164 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4614
timestamp 1711653199
transform 1 0 156 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4615
timestamp 1711653199
transform 1 0 140 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4616
timestamp 1711653199
transform 1 0 140 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4617
timestamp 1711653199
transform 1 0 108 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4618
timestamp 1711653199
transform 1 0 92 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4619
timestamp 1711653199
transform 1 0 380 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4620
timestamp 1711653199
transform 1 0 84 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4621
timestamp 1711653199
transform 1 0 188 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4622
timestamp 1711653199
transform 1 0 132 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_4623
timestamp 1711653199
transform 1 0 196 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4624
timestamp 1711653199
transform 1 0 180 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_4625
timestamp 1711653199
transform 1 0 2972 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4626
timestamp 1711653199
transform 1 0 2924 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4627
timestamp 1711653199
transform 1 0 2500 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_4628
timestamp 1711653199
transform 1 0 1844 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4629
timestamp 1711653199
transform 1 0 1508 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4630
timestamp 1711653199
transform 1 0 916 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4631
timestamp 1711653199
transform 1 0 500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4632
timestamp 1711653199
transform 1 0 284 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4633
timestamp 1711653199
transform 1 0 212 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4634
timestamp 1711653199
transform 1 0 756 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4635
timestamp 1711653199
transform 1 0 388 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4636
timestamp 1711653199
transform 1 0 2324 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4637
timestamp 1711653199
transform 1 0 2300 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4638
timestamp 1711653199
transform 1 0 2220 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4639
timestamp 1711653199
transform 1 0 2148 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_4640
timestamp 1711653199
transform 1 0 1684 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4641
timestamp 1711653199
transform 1 0 1292 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4642
timestamp 1711653199
transform 1 0 876 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4643
timestamp 1711653199
transform 1 0 124 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4644
timestamp 1711653199
transform 1 0 124 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4645
timestamp 1711653199
transform 1 0 124 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4646
timestamp 1711653199
transform 1 0 92 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4647
timestamp 1711653199
transform 1 0 92 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4648
timestamp 1711653199
transform 1 0 84 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4649
timestamp 1711653199
transform 1 0 356 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4650
timestamp 1711653199
transform 1 0 84 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4651
timestamp 1711653199
transform 1 0 164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4652
timestamp 1711653199
transform 1 0 124 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4653
timestamp 1711653199
transform 1 0 404 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4654
timestamp 1711653199
transform 1 0 388 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4655
timestamp 1711653199
transform 1 0 356 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4656
timestamp 1711653199
transform 1 0 820 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4657
timestamp 1711653199
transform 1 0 396 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4658
timestamp 1711653199
transform 1 0 1460 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4659
timestamp 1711653199
transform 1 0 836 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4660
timestamp 1711653199
transform 1 0 740 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4661
timestamp 1711653199
transform 1 0 684 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4662
timestamp 1711653199
transform 1 0 596 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4663
timestamp 1711653199
transform 1 0 540 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4664
timestamp 1711653199
transform 1 0 452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4665
timestamp 1711653199
transform 1 0 460 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4666
timestamp 1711653199
transform 1 0 460 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4667
timestamp 1711653199
transform 1 0 476 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4668
timestamp 1711653199
transform 1 0 444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4669
timestamp 1711653199
transform 1 0 572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4670
timestamp 1711653199
transform 1 0 404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4671
timestamp 1711653199
transform 1 0 396 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4672
timestamp 1711653199
transform 1 0 348 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4673
timestamp 1711653199
transform 1 0 348 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4674
timestamp 1711653199
transform 1 0 212 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4675
timestamp 1711653199
transform 1 0 132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4676
timestamp 1711653199
transform 1 0 236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4677
timestamp 1711653199
transform 1 0 188 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4678
timestamp 1711653199
transform 1 0 476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4679
timestamp 1711653199
transform 1 0 460 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4680
timestamp 1711653199
transform 1 0 316 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4681
timestamp 1711653199
transform 1 0 292 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_4682
timestamp 1711653199
transform 1 0 292 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4683
timestamp 1711653199
transform 1 0 476 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4684
timestamp 1711653199
transform 1 0 452 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4685
timestamp 1711653199
transform 1 0 924 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4686
timestamp 1711653199
transform 1 0 460 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4687
timestamp 1711653199
transform 1 0 1540 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4688
timestamp 1711653199
transform 1 0 1540 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4689
timestamp 1711653199
transform 1 0 1436 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_4690
timestamp 1711653199
transform 1 0 788 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4691
timestamp 1711653199
transform 1 0 396 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4692
timestamp 1711653199
transform 1 0 396 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4693
timestamp 1711653199
transform 1 0 2068 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4694
timestamp 1711653199
transform 1 0 1668 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4695
timestamp 1711653199
transform 1 0 1452 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4696
timestamp 1711653199
transform 1 0 908 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4697
timestamp 1711653199
transform 1 0 956 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4698
timestamp 1711653199
transform 1 0 876 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_4699
timestamp 1711653199
transform 1 0 2404 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4700
timestamp 1711653199
transform 1 0 2380 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4701
timestamp 1711653199
transform 1 0 2084 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4702
timestamp 1711653199
transform 1 0 2084 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_4703
timestamp 1711653199
transform 1 0 1740 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4704
timestamp 1711653199
transform 1 0 1700 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4705
timestamp 1711653199
transform 1 0 1268 0 1 2085
box -2 -2 2 2
use M2_M1  M2_M1_4706
timestamp 1711653199
transform 1 0 1268 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4707
timestamp 1711653199
transform 1 0 2116 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4708
timestamp 1711653199
transform 1 0 1964 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_4709
timestamp 1711653199
transform 1 0 1044 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4710
timestamp 1711653199
transform 1 0 868 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4711
timestamp 1711653199
transform 1 0 572 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4712
timestamp 1711653199
transform 1 0 548 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4713
timestamp 1711653199
transform 1 0 484 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_4714
timestamp 1711653199
transform 1 0 556 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4715
timestamp 1711653199
transform 1 0 524 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4716
timestamp 1711653199
transform 1 0 772 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4717
timestamp 1711653199
transform 1 0 516 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4718
timestamp 1711653199
transform 1 0 540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4719
timestamp 1711653199
transform 1 0 524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4720
timestamp 1711653199
transform 1 0 620 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4721
timestamp 1711653199
transform 1 0 580 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4722
timestamp 1711653199
transform 1 0 596 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_4723
timestamp 1711653199
transform 1 0 468 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4724
timestamp 1711653199
transform 1 0 1036 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4725
timestamp 1711653199
transform 1 0 876 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4726
timestamp 1711653199
transform 1 0 564 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4727
timestamp 1711653199
transform 1 0 524 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4728
timestamp 1711653199
transform 1 0 500 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4729
timestamp 1711653199
transform 1 0 924 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_4730
timestamp 1711653199
transform 1 0 868 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4731
timestamp 1711653199
transform 1 0 748 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4732
timestamp 1711653199
transform 1 0 668 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4733
timestamp 1711653199
transform 1 0 740 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4734
timestamp 1711653199
transform 1 0 676 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_4735
timestamp 1711653199
transform 1 0 708 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4736
timestamp 1711653199
transform 1 0 708 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4737
timestamp 1711653199
transform 1 0 836 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4738
timestamp 1711653199
transform 1 0 740 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4739
timestamp 1711653199
transform 1 0 844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_4740
timestamp 1711653199
transform 1 0 724 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4741
timestamp 1711653199
transform 1 0 916 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4742
timestamp 1711653199
transform 1 0 884 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4743
timestamp 1711653199
transform 1 0 524 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4744
timestamp 1711653199
transform 1 0 516 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4745
timestamp 1711653199
transform 1 0 1108 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4746
timestamp 1711653199
transform 1 0 996 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4747
timestamp 1711653199
transform 1 0 1100 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4748
timestamp 1711653199
transform 1 0 1068 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4749
timestamp 1711653199
transform 1 0 2372 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4750
timestamp 1711653199
transform 1 0 2268 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4751
timestamp 1711653199
transform 1 0 2220 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4752
timestamp 1711653199
transform 1 0 2004 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4753
timestamp 1711653199
transform 1 0 1828 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4754
timestamp 1711653199
transform 1 0 1228 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_4755
timestamp 1711653199
transform 1 0 1180 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_4756
timestamp 1711653199
transform 1 0 1180 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4757
timestamp 1711653199
transform 1 0 444 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4758
timestamp 1711653199
transform 1 0 436 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4759
timestamp 1711653199
transform 1 0 484 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4760
timestamp 1711653199
transform 1 0 412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4761
timestamp 1711653199
transform 1 0 516 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4762
timestamp 1711653199
transform 1 0 388 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4763
timestamp 1711653199
transform 1 0 420 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4764
timestamp 1711653199
transform 1 0 404 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4765
timestamp 1711653199
transform 1 0 852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4766
timestamp 1711653199
transform 1 0 652 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_4767
timestamp 1711653199
transform 1 0 468 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4768
timestamp 1711653199
transform 1 0 852 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_4769
timestamp 1711653199
transform 1 0 716 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4770
timestamp 1711653199
transform 1 0 700 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4771
timestamp 1711653199
transform 1 0 492 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_4772
timestamp 1711653199
transform 1 0 436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4773
timestamp 1711653199
transform 1 0 724 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_4774
timestamp 1711653199
transform 1 0 692 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4775
timestamp 1711653199
transform 1 0 548 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4776
timestamp 1711653199
transform 1 0 548 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_4777
timestamp 1711653199
transform 1 0 540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4778
timestamp 1711653199
transform 1 0 540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4779
timestamp 1711653199
transform 1 0 628 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4780
timestamp 1711653199
transform 1 0 628 0 1 1685
box -2 -2 2 2
use M2_M1  M2_M1_4781
timestamp 1711653199
transform 1 0 596 0 1 1685
box -2 -2 2 2
use M2_M1  M2_M1_4782
timestamp 1711653199
transform 1 0 564 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_4783
timestamp 1711653199
transform 1 0 628 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4784
timestamp 1711653199
transform 1 0 580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4785
timestamp 1711653199
transform 1 0 516 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4786
timestamp 1711653199
transform 1 0 444 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4787
timestamp 1711653199
transform 1 0 724 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4788
timestamp 1711653199
transform 1 0 436 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4789
timestamp 1711653199
transform 1 0 596 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_4790
timestamp 1711653199
transform 1 0 556 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_4791
timestamp 1711653199
transform 1 0 804 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4792
timestamp 1711653199
transform 1 0 716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4793
timestamp 1711653199
transform 1 0 684 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4794
timestamp 1711653199
transform 1 0 636 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4795
timestamp 1711653199
transform 1 0 612 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4796
timestamp 1711653199
transform 1 0 556 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4797
timestamp 1711653199
transform 1 0 516 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4798
timestamp 1711653199
transform 1 0 628 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_4799
timestamp 1711653199
transform 1 0 492 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4800
timestamp 1711653199
transform 1 0 516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4801
timestamp 1711653199
transform 1 0 500 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_4802
timestamp 1711653199
transform 1 0 700 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4803
timestamp 1711653199
transform 1 0 524 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4804
timestamp 1711653199
transform 1 0 572 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4805
timestamp 1711653199
transform 1 0 564 0 1 1285
box -2 -2 2 2
use M2_M1  M2_M1_4806
timestamp 1711653199
transform 1 0 900 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4807
timestamp 1711653199
transform 1 0 844 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4808
timestamp 1711653199
transform 1 0 812 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4809
timestamp 1711653199
transform 1 0 1060 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_4810
timestamp 1711653199
transform 1 0 1004 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4811
timestamp 1711653199
transform 1 0 684 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4812
timestamp 1711653199
transform 1 0 636 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_4813
timestamp 1711653199
transform 1 0 636 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_4814
timestamp 1711653199
transform 1 0 1764 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4815
timestamp 1711653199
transform 1 0 1052 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4816
timestamp 1711653199
transform 1 0 988 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4817
timestamp 1711653199
transform 1 0 964 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4818
timestamp 1711653199
transform 1 0 964 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_4819
timestamp 1711653199
transform 1 0 932 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4820
timestamp 1711653199
transform 1 0 924 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_4821
timestamp 1711653199
transform 1 0 948 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4822
timestamp 1711653199
transform 1 0 932 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_4823
timestamp 1711653199
transform 1 0 940 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4824
timestamp 1711653199
transform 1 0 940 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4825
timestamp 1711653199
transform 1 0 772 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4826
timestamp 1711653199
transform 1 0 612 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4827
timestamp 1711653199
transform 1 0 612 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4828
timestamp 1711653199
transform 1 0 596 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_4829
timestamp 1711653199
transform 1 0 1204 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4830
timestamp 1711653199
transform 1 0 628 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4831
timestamp 1711653199
transform 1 0 532 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4832
timestamp 1711653199
transform 1 0 484 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4833
timestamp 1711653199
transform 1 0 1780 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4834
timestamp 1711653199
transform 1 0 1380 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_4835
timestamp 1711653199
transform 1 0 1332 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4836
timestamp 1711653199
transform 1 0 980 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4837
timestamp 1711653199
transform 1 0 1756 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4838
timestamp 1711653199
transform 1 0 1740 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4839
timestamp 1711653199
transform 1 0 1748 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4840
timestamp 1711653199
transform 1 0 1748 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4841
timestamp 1711653199
transform 1 0 1740 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_4842
timestamp 1711653199
transform 1 0 1716 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_4843
timestamp 1711653199
transform 1 0 2268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4844
timestamp 1711653199
transform 1 0 1844 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4845
timestamp 1711653199
transform 1 0 2108 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_4846
timestamp 1711653199
transform 1 0 2100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4847
timestamp 1711653199
transform 1 0 1852 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4848
timestamp 1711653199
transform 1 0 1756 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4849
timestamp 1711653199
transform 1 0 1748 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4850
timestamp 1711653199
transform 1 0 1732 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4851
timestamp 1711653199
transform 1 0 1460 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_4852
timestamp 1711653199
transform 1 0 1412 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4853
timestamp 1711653199
transform 1 0 1420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4854
timestamp 1711653199
transform 1 0 1404 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_4855
timestamp 1711653199
transform 1 0 2188 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4856
timestamp 1711653199
transform 1 0 1756 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4857
timestamp 1711653199
transform 1 0 1820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4858
timestamp 1711653199
transform 1 0 1820 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4859
timestamp 1711653199
transform 1 0 2220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_4860
timestamp 1711653199
transform 1 0 2220 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_4861
timestamp 1711653199
transform 1 0 1652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4862
timestamp 1711653199
transform 1 0 1548 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4863
timestamp 1711653199
transform 1 0 1588 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4864
timestamp 1711653199
transform 1 0 1580 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_4865
timestamp 1711653199
transform 1 0 1332 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4866
timestamp 1711653199
transform 1 0 1164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4867
timestamp 1711653199
transform 1 0 932 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4868
timestamp 1711653199
transform 1 0 1980 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4869
timestamp 1711653199
transform 1 0 1732 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4870
timestamp 1711653199
transform 1 0 1404 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4871
timestamp 1711653199
transform 1 0 1372 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_4872
timestamp 1711653199
transform 1 0 1164 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4873
timestamp 1711653199
transform 1 0 964 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4874
timestamp 1711653199
transform 1 0 644 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4875
timestamp 1711653199
transform 1 0 628 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4876
timestamp 1711653199
transform 1 0 1644 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4877
timestamp 1711653199
transform 1 0 788 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4878
timestamp 1711653199
transform 1 0 948 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4879
timestamp 1711653199
transform 1 0 924 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4880
timestamp 1711653199
transform 1 0 860 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4881
timestamp 1711653199
transform 1 0 796 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_4882
timestamp 1711653199
transform 1 0 804 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4883
timestamp 1711653199
transform 1 0 780 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4884
timestamp 1711653199
transform 1 0 844 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4885
timestamp 1711653199
transform 1 0 804 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_4886
timestamp 1711653199
transform 1 0 796 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_4887
timestamp 1711653199
transform 1 0 796 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_4888
timestamp 1711653199
transform 1 0 868 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_4889
timestamp 1711653199
transform 1 0 852 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4890
timestamp 1711653199
transform 1 0 852 0 1 1485
box -2 -2 2 2
use M2_M1  M2_M1_4891
timestamp 1711653199
transform 1 0 852 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4892
timestamp 1711653199
transform 1 0 852 0 1 895
box -2 -2 2 2
use M2_M1  M2_M1_4893
timestamp 1711653199
transform 1 0 852 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_4894
timestamp 1711653199
transform 1 0 836 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_4895
timestamp 1711653199
transform 1 0 828 0 1 1485
box -2 -2 2 2
use M2_M1  M2_M1_4896
timestamp 1711653199
transform 1 0 828 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4897
timestamp 1711653199
transform 1 0 780 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4898
timestamp 1711653199
transform 1 0 772 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4899
timestamp 1711653199
transform 1 0 756 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4900
timestamp 1711653199
transform 1 0 852 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4901
timestamp 1711653199
transform 1 0 852 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4902
timestamp 1711653199
transform 1 0 956 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4903
timestamp 1711653199
transform 1 0 860 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4904
timestamp 1711653199
transform 1 0 852 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4905
timestamp 1711653199
transform 1 0 804 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4906
timestamp 1711653199
transform 1 0 804 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_4907
timestamp 1711653199
transform 1 0 748 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4908
timestamp 1711653199
transform 1 0 748 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4909
timestamp 1711653199
transform 1 0 812 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4910
timestamp 1711653199
transform 1 0 772 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_4911
timestamp 1711653199
transform 1 0 1556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_4912
timestamp 1711653199
transform 1 0 836 0 1 785
box -2 -2 2 2
use M2_M1  M2_M1_4913
timestamp 1711653199
transform 1 0 820 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_4914
timestamp 1711653199
transform 1 0 820 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_4915
timestamp 1711653199
transform 1 0 820 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4916
timestamp 1711653199
transform 1 0 788 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4917
timestamp 1711653199
transform 1 0 516 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4918
timestamp 1711653199
transform 1 0 876 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4919
timestamp 1711653199
transform 1 0 796 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4920
timestamp 1711653199
transform 1 0 812 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4921
timestamp 1711653199
transform 1 0 764 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4922
timestamp 1711653199
transform 1 0 836 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_4923
timestamp 1711653199
transform 1 0 820 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4924
timestamp 1711653199
transform 1 0 820 0 1 1045
box -2 -2 2 2
use M2_M1  M2_M1_4925
timestamp 1711653199
transform 1 0 820 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_4926
timestamp 1711653199
transform 1 0 820 0 1 985
box -2 -2 2 2
use M2_M1  M2_M1_4927
timestamp 1711653199
transform 1 0 804 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_4928
timestamp 1711653199
transform 1 0 772 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4929
timestamp 1711653199
transform 1 0 772 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_4930
timestamp 1711653199
transform 1 0 804 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4931
timestamp 1711653199
transform 1 0 780 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4932
timestamp 1711653199
transform 1 0 828 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4933
timestamp 1711653199
transform 1 0 788 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4934
timestamp 1711653199
transform 1 0 868 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4935
timestamp 1711653199
transform 1 0 748 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_4936
timestamp 1711653199
transform 1 0 804 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_4937
timestamp 1711653199
transform 1 0 772 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4938
timestamp 1711653199
transform 1 0 652 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4939
timestamp 1711653199
transform 1 0 500 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4940
timestamp 1711653199
transform 1 0 436 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4941
timestamp 1711653199
transform 1 0 436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4942
timestamp 1711653199
transform 1 0 388 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4943
timestamp 1711653199
transform 1 0 364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_4944
timestamp 1711653199
transform 1 0 428 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_4945
timestamp 1711653199
transform 1 0 372 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4946
timestamp 1711653199
transform 1 0 444 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_4947
timestamp 1711653199
transform 1 0 436 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4948
timestamp 1711653199
transform 1 0 500 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4949
timestamp 1711653199
transform 1 0 492 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4950
timestamp 1711653199
transform 1 0 428 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_4951
timestamp 1711653199
transform 1 0 388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_4952
timestamp 1711653199
transform 1 0 444 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4953
timestamp 1711653199
transform 1 0 412 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_4954
timestamp 1711653199
transform 1 0 436 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_4955
timestamp 1711653199
transform 1 0 380 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_4956
timestamp 1711653199
transform 1 0 428 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4957
timestamp 1711653199
transform 1 0 420 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4958
timestamp 1711653199
transform 1 0 380 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4959
timestamp 1711653199
transform 1 0 364 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_4960
timestamp 1711653199
transform 1 0 404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4961
timestamp 1711653199
transform 1 0 380 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_4962
timestamp 1711653199
transform 1 0 364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4963
timestamp 1711653199
transform 1 0 300 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_4964
timestamp 1711653199
transform 1 0 212 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_4965
timestamp 1711653199
transform 1 0 372 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_4966
timestamp 1711653199
transform 1 0 356 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_4967
timestamp 1711653199
transform 1 0 452 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4968
timestamp 1711653199
transform 1 0 444 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_4969
timestamp 1711653199
transform 1 0 508 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4970
timestamp 1711653199
transform 1 0 460 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_4971
timestamp 1711653199
transform 1 0 444 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_4972
timestamp 1711653199
transform 1 0 548 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4973
timestamp 1711653199
transform 1 0 484 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4974
timestamp 1711653199
transform 1 0 516 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4975
timestamp 1711653199
transform 1 0 476 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4976
timestamp 1711653199
transform 1 0 428 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_4977
timestamp 1711653199
transform 1 0 404 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_4978
timestamp 1711653199
transform 1 0 844 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4979
timestamp 1711653199
transform 1 0 828 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4980
timestamp 1711653199
transform 1 0 812 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4981
timestamp 1711653199
transform 1 0 716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_4982
timestamp 1711653199
transform 1 0 668 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4983
timestamp 1711653199
transform 1 0 564 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_4984
timestamp 1711653199
transform 1 0 588 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4985
timestamp 1711653199
transform 1 0 180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4986
timestamp 1711653199
transform 1 0 124 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_4987
timestamp 1711653199
transform 1 0 84 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_4988
timestamp 1711653199
transform 1 0 228 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4989
timestamp 1711653199
transform 1 0 148 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4990
timestamp 1711653199
transform 1 0 308 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_4991
timestamp 1711653199
transform 1 0 228 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_4992
timestamp 1711653199
transform 1 0 252 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_4993
timestamp 1711653199
transform 1 0 220 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_4994
timestamp 1711653199
transform 1 0 380 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_4995
timestamp 1711653199
transform 1 0 292 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4996
timestamp 1711653199
transform 1 0 260 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_4997
timestamp 1711653199
transform 1 0 196 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4998
timestamp 1711653199
transform 1 0 148 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_4999
timestamp 1711653199
transform 1 0 340 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5000
timestamp 1711653199
transform 1 0 284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5001
timestamp 1711653199
transform 1 0 284 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5002
timestamp 1711653199
transform 1 0 268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5003
timestamp 1711653199
transform 1 0 364 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5004
timestamp 1711653199
transform 1 0 340 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5005
timestamp 1711653199
transform 1 0 308 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5006
timestamp 1711653199
transform 1 0 300 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5007
timestamp 1711653199
transform 1 0 388 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_5008
timestamp 1711653199
transform 1 0 372 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5009
timestamp 1711653199
transform 1 0 324 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5010
timestamp 1711653199
transform 1 0 316 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5011
timestamp 1711653199
transform 1 0 1332 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5012
timestamp 1711653199
transform 1 0 324 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5013
timestamp 1711653199
transform 1 0 300 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5014
timestamp 1711653199
transform 1 0 196 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5015
timestamp 1711653199
transform 1 0 116 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5016
timestamp 1711653199
transform 1 0 116 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5017
timestamp 1711653199
transform 1 0 196 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5018
timestamp 1711653199
transform 1 0 172 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5019
timestamp 1711653199
transform 1 0 3004 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5020
timestamp 1711653199
transform 1 0 1380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5021
timestamp 1711653199
transform 1 0 1364 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5022
timestamp 1711653199
transform 1 0 284 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5023
timestamp 1711653199
transform 1 0 252 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5024
timestamp 1711653199
transform 1 0 244 0 1 1245
box -2 -2 2 2
use M2_M1  M2_M1_5025
timestamp 1711653199
transform 1 0 228 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5026
timestamp 1711653199
transform 1 0 220 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_5027
timestamp 1711653199
transform 1 0 212 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5028
timestamp 1711653199
transform 1 0 380 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5029
timestamp 1711653199
transform 1 0 260 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5030
timestamp 1711653199
transform 1 0 292 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5031
timestamp 1711653199
transform 1 0 284 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5032
timestamp 1711653199
transform 1 0 268 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_5033
timestamp 1711653199
transform 1 0 260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5034
timestamp 1711653199
transform 1 0 1036 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5035
timestamp 1711653199
transform 1 0 692 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5036
timestamp 1711653199
transform 1 0 596 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5037
timestamp 1711653199
transform 1 0 668 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5038
timestamp 1711653199
transform 1 0 388 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5039
timestamp 1711653199
transform 1 0 1452 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5040
timestamp 1711653199
transform 1 0 1444 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5041
timestamp 1711653199
transform 1 0 1396 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5042
timestamp 1711653199
transform 1 0 1388 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5043
timestamp 1711653199
transform 1 0 1412 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5044
timestamp 1711653199
transform 1 0 1348 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5045
timestamp 1711653199
transform 1 0 1388 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5046
timestamp 1711653199
transform 1 0 1364 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5047
timestamp 1711653199
transform 1 0 1396 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5048
timestamp 1711653199
transform 1 0 1276 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5049
timestamp 1711653199
transform 1 0 1252 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5050
timestamp 1711653199
transform 1 0 1388 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5051
timestamp 1711653199
transform 1 0 1388 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5052
timestamp 1711653199
transform 1 0 2412 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5053
timestamp 1711653199
transform 1 0 2396 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5054
timestamp 1711653199
transform 1 0 2300 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5055
timestamp 1711653199
transform 1 0 2204 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5056
timestamp 1711653199
transform 1 0 1404 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5057
timestamp 1711653199
transform 1 0 1340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5058
timestamp 1711653199
transform 1 0 1316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5059
timestamp 1711653199
transform 1 0 1300 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5060
timestamp 1711653199
transform 1 0 1396 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5061
timestamp 1711653199
transform 1 0 1380 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5062
timestamp 1711653199
transform 1 0 1420 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5063
timestamp 1711653199
transform 1 0 1404 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5064
timestamp 1711653199
transform 1 0 1444 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5065
timestamp 1711653199
transform 1 0 1428 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5066
timestamp 1711653199
transform 1 0 1404 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5067
timestamp 1711653199
transform 1 0 1404 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5068
timestamp 1711653199
transform 1 0 1364 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5069
timestamp 1711653199
transform 1 0 1364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5070
timestamp 1711653199
transform 1 0 1372 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5071
timestamp 1711653199
transform 1 0 1348 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5072
timestamp 1711653199
transform 1 0 1412 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5073
timestamp 1711653199
transform 1 0 1340 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5074
timestamp 1711653199
transform 1 0 1476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5075
timestamp 1711653199
transform 1 0 1380 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5076
timestamp 1711653199
transform 1 0 1316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5077
timestamp 1711653199
transform 1 0 1252 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5078
timestamp 1711653199
transform 1 0 1164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5079
timestamp 1711653199
transform 1 0 1476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5080
timestamp 1711653199
transform 1 0 1444 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5081
timestamp 1711653199
transform 1 0 1460 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5082
timestamp 1711653199
transform 1 0 1460 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5083
timestamp 1711653199
transform 1 0 2476 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5084
timestamp 1711653199
transform 1 0 2396 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5085
timestamp 1711653199
transform 1 0 2228 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5086
timestamp 1711653199
transform 1 0 2212 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5087
timestamp 1711653199
transform 1 0 1500 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5088
timestamp 1711653199
transform 1 0 1460 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5089
timestamp 1711653199
transform 1 0 1388 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5090
timestamp 1711653199
transform 1 0 1188 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5091
timestamp 1711653199
transform 1 0 2044 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5092
timestamp 1711653199
transform 1 0 2044 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5093
timestamp 1711653199
transform 1 0 2012 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5094
timestamp 1711653199
transform 1 0 1516 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5095
timestamp 1711653199
transform 1 0 1476 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5096
timestamp 1711653199
transform 1 0 1268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5097
timestamp 1711653199
transform 1 0 1340 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5098
timestamp 1711653199
transform 1 0 1180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5099
timestamp 1711653199
transform 1 0 1156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5100
timestamp 1711653199
transform 1 0 1148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5101
timestamp 1711653199
transform 1 0 1140 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5102
timestamp 1711653199
transform 1 0 1140 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5103
timestamp 1711653199
transform 1 0 1052 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5104
timestamp 1711653199
transform 1 0 956 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5105
timestamp 1711653199
transform 1 0 1108 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5106
timestamp 1711653199
transform 1 0 1100 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5107
timestamp 1711653199
transform 1 0 1340 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5108
timestamp 1711653199
transform 1 0 1332 0 1 1955
box -2 -2 2 2
use M2_M1  M2_M1_5109
timestamp 1711653199
transform 1 0 1252 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5110
timestamp 1711653199
transform 1 0 1188 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5111
timestamp 1711653199
transform 1 0 1164 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5112
timestamp 1711653199
transform 1 0 1228 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5113
timestamp 1711653199
transform 1 0 1172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5114
timestamp 1711653199
transform 1 0 1124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5115
timestamp 1711653199
transform 1 0 1036 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5116
timestamp 1711653199
transform 1 0 996 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5117
timestamp 1711653199
transform 1 0 980 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5118
timestamp 1711653199
transform 1 0 996 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5119
timestamp 1711653199
transform 1 0 996 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_5120
timestamp 1711653199
transform 1 0 988 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5121
timestamp 1711653199
transform 1 0 988 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5122
timestamp 1711653199
transform 1 0 1252 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5123
timestamp 1711653199
transform 1 0 1124 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5124
timestamp 1711653199
transform 1 0 1084 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5125
timestamp 1711653199
transform 1 0 996 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5126
timestamp 1711653199
transform 1 0 964 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5127
timestamp 1711653199
transform 1 0 964 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5128
timestamp 1711653199
transform 1 0 940 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5129
timestamp 1711653199
transform 1 0 940 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5130
timestamp 1711653199
transform 1 0 1212 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5131
timestamp 1711653199
transform 1 0 1148 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5132
timestamp 1711653199
transform 1 0 1332 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5133
timestamp 1711653199
transform 1 0 1276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5134
timestamp 1711653199
transform 1 0 1316 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5135
timestamp 1711653199
transform 1 0 1276 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5136
timestamp 1711653199
transform 1 0 1860 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5137
timestamp 1711653199
transform 1 0 1516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5138
timestamp 1711653199
transform 1 0 1956 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5139
timestamp 1711653199
transform 1 0 1852 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5140
timestamp 1711653199
transform 1 0 2892 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5141
timestamp 1711653199
transform 1 0 2860 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5142
timestamp 1711653199
transform 1 0 2764 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5143
timestamp 1711653199
transform 1 0 2668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5144
timestamp 1711653199
transform 1 0 2612 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5145
timestamp 1711653199
transform 1 0 2324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5146
timestamp 1711653199
transform 1 0 2148 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5147
timestamp 1711653199
transform 1 0 1956 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5148
timestamp 1711653199
transform 1 0 1940 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5149
timestamp 1711653199
transform 1 0 1652 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5150
timestamp 1711653199
transform 1 0 1372 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5151
timestamp 1711653199
transform 1 0 1348 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5152
timestamp 1711653199
transform 1 0 1308 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5153
timestamp 1711653199
transform 1 0 1316 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5154
timestamp 1711653199
transform 1 0 1316 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5155
timestamp 1711653199
transform 1 0 1260 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5156
timestamp 1711653199
transform 1 0 1244 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5157
timestamp 1711653199
transform 1 0 1324 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5158
timestamp 1711653199
transform 1 0 1316 0 1 1255
box -2 -2 2 2
use M2_M1  M2_M1_5159
timestamp 1711653199
transform 1 0 1300 0 1 1255
box -2 -2 2 2
use M2_M1  M2_M1_5160
timestamp 1711653199
transform 1 0 1300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5161
timestamp 1711653199
transform 1 0 1332 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5162
timestamp 1711653199
transform 1 0 1276 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5163
timestamp 1711653199
transform 1 0 1236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5164
timestamp 1711653199
transform 1 0 1260 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5165
timestamp 1711653199
transform 1 0 1244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5166
timestamp 1711653199
transform 1 0 1236 0 1 855
box -2 -2 2 2
use M2_M1  M2_M1_5167
timestamp 1711653199
transform 1 0 1212 0 1 855
box -2 -2 2 2
use M2_M1  M2_M1_5168
timestamp 1711653199
transform 1 0 1212 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5169
timestamp 1711653199
transform 1 0 1116 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5170
timestamp 1711653199
transform 1 0 1116 0 1 505
box -2 -2 2 2
use M2_M1  M2_M1_5171
timestamp 1711653199
transform 1 0 1148 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5172
timestamp 1711653199
transform 1 0 1148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5173
timestamp 1711653199
transform 1 0 1140 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5174
timestamp 1711653199
transform 1 0 1132 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5175
timestamp 1711653199
transform 1 0 1220 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5176
timestamp 1711653199
transform 1 0 1140 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_5177
timestamp 1711653199
transform 1 0 1236 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5178
timestamp 1711653199
transform 1 0 1236 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5179
timestamp 1711653199
transform 1 0 1276 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_5180
timestamp 1711653199
transform 1 0 1268 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5181
timestamp 1711653199
transform 1 0 1300 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5182
timestamp 1711653199
transform 1 0 1292 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5183
timestamp 1711653199
transform 1 0 1236 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5184
timestamp 1711653199
transform 1 0 1236 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5185
timestamp 1711653199
transform 1 0 2996 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5186
timestamp 1711653199
transform 1 0 2860 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5187
timestamp 1711653199
transform 1 0 2420 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5188
timestamp 1711653199
transform 1 0 2180 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5189
timestamp 1711653199
transform 1 0 1420 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5190
timestamp 1711653199
transform 1 0 1764 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5191
timestamp 1711653199
transform 1 0 1700 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5192
timestamp 1711653199
transform 1 0 2380 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5193
timestamp 1711653199
transform 1 0 2116 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5194
timestamp 1711653199
transform 1 0 1724 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5195
timestamp 1711653199
transform 1 0 1788 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5196
timestamp 1711653199
transform 1 0 1764 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5197
timestamp 1711653199
transform 1 0 1412 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5198
timestamp 1711653199
transform 1 0 1116 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5199
timestamp 1711653199
transform 1 0 1084 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_5200
timestamp 1711653199
transform 1 0 1076 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5201
timestamp 1711653199
transform 1 0 1012 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5202
timestamp 1711653199
transform 1 0 1012 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5203
timestamp 1711653199
transform 1 0 1060 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5204
timestamp 1711653199
transform 1 0 1052 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5205
timestamp 1711653199
transform 1 0 1164 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5206
timestamp 1711653199
transform 1 0 1132 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5207
timestamp 1711653199
transform 1 0 1116 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5208
timestamp 1711653199
transform 1 0 1020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5209
timestamp 1711653199
transform 1 0 1156 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_5210
timestamp 1711653199
transform 1 0 1124 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_5211
timestamp 1711653199
transform 1 0 1124 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5212
timestamp 1711653199
transform 1 0 1100 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5213
timestamp 1711653199
transform 1 0 1068 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5214
timestamp 1711653199
transform 1 0 1060 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5215
timestamp 1711653199
transform 1 0 980 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5216
timestamp 1711653199
transform 1 0 1964 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5217
timestamp 1711653199
transform 1 0 1612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5218
timestamp 1711653199
transform 1 0 1092 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5219
timestamp 1711653199
transform 1 0 1092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5220
timestamp 1711653199
transform 1 0 1108 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5221
timestamp 1711653199
transform 1 0 1100 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_5222
timestamp 1711653199
transform 1 0 1180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5223
timestamp 1711653199
transform 1 0 1156 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5224
timestamp 1711653199
transform 1 0 1060 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_5225
timestamp 1711653199
transform 1 0 1060 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5226
timestamp 1711653199
transform 1 0 1044 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5227
timestamp 1711653199
transform 1 0 956 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5228
timestamp 1711653199
transform 1 0 1116 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5229
timestamp 1711653199
transform 1 0 1068 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5230
timestamp 1711653199
transform 1 0 2484 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5231
timestamp 1711653199
transform 1 0 2356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5232
timestamp 1711653199
transform 1 0 2092 0 1 1924
box -2 -2 2 2
use M2_M1  M2_M1_5233
timestamp 1711653199
transform 1 0 1348 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5234
timestamp 1711653199
transform 1 0 1844 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5235
timestamp 1711653199
transform 1 0 1780 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5236
timestamp 1711653199
transform 1 0 2148 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5237
timestamp 1711653199
transform 1 0 2044 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5238
timestamp 1711653199
transform 1 0 1812 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5239
timestamp 1711653199
transform 1 0 1876 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5240
timestamp 1711653199
transform 1 0 1852 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_5241
timestamp 1711653199
transform 1 0 2436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5242
timestamp 1711653199
transform 1 0 2268 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5243
timestamp 1711653199
transform 1 0 2404 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5244
timestamp 1711653199
transform 1 0 2404 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5245
timestamp 1711653199
transform 1 0 2532 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5246
timestamp 1711653199
transform 1 0 2412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5247
timestamp 1711653199
transform 1 0 2548 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5248
timestamp 1711653199
transform 1 0 2540 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5249
timestamp 1711653199
transform 1 0 2564 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5250
timestamp 1711653199
transform 1 0 2492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5251
timestamp 1711653199
transform 1 0 2316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5252
timestamp 1711653199
transform 1 0 2268 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5253
timestamp 1711653199
transform 1 0 2252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_5254
timestamp 1711653199
transform 1 0 2052 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5255
timestamp 1711653199
transform 1 0 1956 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5256
timestamp 1711653199
transform 1 0 2604 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_5257
timestamp 1711653199
transform 1 0 2548 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5258
timestamp 1711653199
transform 1 0 2596 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_5259
timestamp 1711653199
transform 1 0 2596 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5260
timestamp 1711653199
transform 1 0 2564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5261
timestamp 1711653199
transform 1 0 2244 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5262
timestamp 1711653199
transform 1 0 2228 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5263
timestamp 1711653199
transform 1 0 2532 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_5264
timestamp 1711653199
transform 1 0 2436 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5265
timestamp 1711653199
transform 1 0 2380 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5266
timestamp 1711653199
transform 1 0 2132 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_5267
timestamp 1711653199
transform 1 0 2348 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_5268
timestamp 1711653199
transform 1 0 2300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5269
timestamp 1711653199
transform 1 0 2236 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5270
timestamp 1711653199
transform 1 0 2196 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5271
timestamp 1711653199
transform 1 0 2692 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5272
timestamp 1711653199
transform 1 0 2636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5273
timestamp 1711653199
transform 1 0 2540 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5274
timestamp 1711653199
transform 1 0 2524 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5275
timestamp 1711653199
transform 1 0 2516 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5276
timestamp 1711653199
transform 1 0 2268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5277
timestamp 1711653199
transform 1 0 2252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5278
timestamp 1711653199
transform 1 0 2012 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5279
timestamp 1711653199
transform 1 0 2028 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5280
timestamp 1711653199
transform 1 0 2028 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5281
timestamp 1711653199
transform 1 0 2036 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5282
timestamp 1711653199
transform 1 0 2036 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5283
timestamp 1711653199
transform 1 0 2868 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5284
timestamp 1711653199
transform 1 0 2868 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5285
timestamp 1711653199
transform 1 0 2828 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5286
timestamp 1711653199
transform 1 0 2828 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5287
timestamp 1711653199
transform 1 0 2788 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5288
timestamp 1711653199
transform 1 0 2676 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_5289
timestamp 1711653199
transform 1 0 2580 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5290
timestamp 1711653199
transform 1 0 2292 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5291
timestamp 1711653199
transform 1 0 2276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5292
timestamp 1711653199
transform 1 0 2276 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5293
timestamp 1711653199
transform 1 0 2012 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5294
timestamp 1711653199
transform 1 0 1596 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5295
timestamp 1711653199
transform 1 0 1980 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5296
timestamp 1711653199
transform 1 0 1932 0 1 2195
box -2 -2 2 2
use M2_M1  M2_M1_5297
timestamp 1711653199
transform 1 0 3116 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5298
timestamp 1711653199
transform 1 0 2316 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5299
timestamp 1711653199
transform 1 0 3044 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5300
timestamp 1711653199
transform 1 0 3036 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5301
timestamp 1711653199
transform 1 0 3196 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5302
timestamp 1711653199
transform 1 0 3052 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5303
timestamp 1711653199
transform 1 0 3188 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5304
timestamp 1711653199
transform 1 0 3148 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5305
timestamp 1711653199
transform 1 0 3148 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5306
timestamp 1711653199
transform 1 0 3140 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5307
timestamp 1711653199
transform 1 0 3180 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_5308
timestamp 1711653199
transform 1 0 3164 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5309
timestamp 1711653199
transform 1 0 3164 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_5310
timestamp 1711653199
transform 1 0 3148 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5311
timestamp 1711653199
transform 1 0 3148 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5312
timestamp 1711653199
transform 1 0 3116 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5313
timestamp 1711653199
transform 1 0 3108 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5314
timestamp 1711653199
transform 1 0 3084 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5315
timestamp 1711653199
transform 1 0 3084 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5316
timestamp 1711653199
transform 1 0 3172 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5317
timestamp 1711653199
transform 1 0 3132 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5318
timestamp 1711653199
transform 1 0 3172 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_5319
timestamp 1711653199
transform 1 0 3060 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5320
timestamp 1711653199
transform 1 0 3044 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5321
timestamp 1711653199
transform 1 0 3044 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5322
timestamp 1711653199
transform 1 0 3044 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5323
timestamp 1711653199
transform 1 0 2956 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5324
timestamp 1711653199
transform 1 0 2556 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5325
timestamp 1711653199
transform 1 0 3204 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5326
timestamp 1711653199
transform 1 0 3196 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5327
timestamp 1711653199
transform 1 0 3212 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5328
timestamp 1711653199
transform 1 0 3124 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5329
timestamp 1711653199
transform 1 0 3140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5330
timestamp 1711653199
transform 1 0 3140 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5331
timestamp 1711653199
transform 1 0 3092 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5332
timestamp 1711653199
transform 1 0 3068 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5333
timestamp 1711653199
transform 1 0 3108 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5334
timestamp 1711653199
transform 1 0 3036 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5335
timestamp 1711653199
transform 1 0 3052 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5336
timestamp 1711653199
transform 1 0 2980 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5337
timestamp 1711653199
transform 1 0 3124 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5338
timestamp 1711653199
transform 1 0 3060 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_5339
timestamp 1711653199
transform 1 0 3004 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5340
timestamp 1711653199
transform 1 0 2948 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5341
timestamp 1711653199
transform 1 0 3156 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5342
timestamp 1711653199
transform 1 0 3076 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5343
timestamp 1711653199
transform 1 0 3132 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5344
timestamp 1711653199
transform 1 0 3044 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5345
timestamp 1711653199
transform 1 0 3156 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5346
timestamp 1711653199
transform 1 0 2460 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5347
timestamp 1711653199
transform 1 0 3396 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_5348
timestamp 1711653199
transform 1 0 3380 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_5349
timestamp 1711653199
transform 1 0 3300 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5350
timestamp 1711653199
transform 1 0 2620 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5351
timestamp 1711653199
transform 1 0 3244 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5352
timestamp 1711653199
transform 1 0 3244 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5353
timestamp 1711653199
transform 1 0 3300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5354
timestamp 1711653199
transform 1 0 3284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5355
timestamp 1711653199
transform 1 0 3316 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_5356
timestamp 1711653199
transform 1 0 3316 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5357
timestamp 1711653199
transform 1 0 3292 0 1 1155
box -2 -2 2 2
use M2_M1  M2_M1_5358
timestamp 1711653199
transform 1 0 3276 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5359
timestamp 1711653199
transform 1 0 3396 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5360
timestamp 1711653199
transform 1 0 3284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5361
timestamp 1711653199
transform 1 0 3340 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5362
timestamp 1711653199
transform 1 0 3324 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5363
timestamp 1711653199
transform 1 0 3284 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5364
timestamp 1711653199
transform 1 0 3284 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_5365
timestamp 1711653199
transform 1 0 3228 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5366
timestamp 1711653199
transform 1 0 3324 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5367
timestamp 1711653199
transform 1 0 3324 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5368
timestamp 1711653199
transform 1 0 3308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5369
timestamp 1711653199
transform 1 0 3308 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5370
timestamp 1711653199
transform 1 0 3324 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5371
timestamp 1711653199
transform 1 0 3308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5372
timestamp 1711653199
transform 1 0 3332 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5373
timestamp 1711653199
transform 1 0 3308 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5374
timestamp 1711653199
transform 1 0 3292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5375
timestamp 1711653199
transform 1 0 3276 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5376
timestamp 1711653199
transform 1 0 3268 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5377
timestamp 1711653199
transform 1 0 3300 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5378
timestamp 1711653199
transform 1 0 3276 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5379
timestamp 1711653199
transform 1 0 3292 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5380
timestamp 1711653199
transform 1 0 3212 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_5381
timestamp 1711653199
transform 1 0 3308 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5382
timestamp 1711653199
transform 1 0 3252 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5383
timestamp 1711653199
transform 1 0 3132 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_5384
timestamp 1711653199
transform 1 0 3188 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5385
timestamp 1711653199
transform 1 0 3164 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5386
timestamp 1711653199
transform 1 0 3252 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5387
timestamp 1711653199
transform 1 0 3252 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5388
timestamp 1711653199
transform 1 0 3268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5389
timestamp 1711653199
transform 1 0 3196 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_5390
timestamp 1711653199
transform 1 0 2932 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5391
timestamp 1711653199
transform 1 0 2932 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5392
timestamp 1711653199
transform 1 0 2820 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5393
timestamp 1711653199
transform 1 0 2572 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5394
timestamp 1711653199
transform 1 0 2380 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5395
timestamp 1711653199
transform 1 0 3164 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5396
timestamp 1711653199
transform 1 0 2372 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5397
timestamp 1711653199
transform 1 0 3172 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5398
timestamp 1711653199
transform 1 0 2676 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_5399
timestamp 1711653199
transform 1 0 3212 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5400
timestamp 1711653199
transform 1 0 3148 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5401
timestamp 1711653199
transform 1 0 3228 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5402
timestamp 1711653199
transform 1 0 3156 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5403
timestamp 1711653199
transform 1 0 3244 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5404
timestamp 1711653199
transform 1 0 3212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5405
timestamp 1711653199
transform 1 0 3260 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5406
timestamp 1711653199
transform 1 0 3260 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_5407
timestamp 1711653199
transform 1 0 3380 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5408
timestamp 1711653199
transform 1 0 3356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5409
timestamp 1711653199
transform 1 0 3348 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5410
timestamp 1711653199
transform 1 0 3348 0 1 1385
box -2 -2 2 2
use M2_M1  M2_M1_5411
timestamp 1711653199
transform 1 0 3348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5412
timestamp 1711653199
transform 1 0 3340 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5413
timestamp 1711653199
transform 1 0 3332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5414
timestamp 1711653199
transform 1 0 3396 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5415
timestamp 1711653199
transform 1 0 3380 0 1 1495
box -2 -2 2 2
use M2_M1  M2_M1_5416
timestamp 1711653199
transform 1 0 3380 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5417
timestamp 1711653199
transform 1 0 3340 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5418
timestamp 1711653199
transform 1 0 3356 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5419
timestamp 1711653199
transform 1 0 3356 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5420
timestamp 1711653199
transform 1 0 3380 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5421
timestamp 1711653199
transform 1 0 3364 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5422
timestamp 1711653199
transform 1 0 3340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5423
timestamp 1711653199
transform 1 0 3252 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5424
timestamp 1711653199
transform 1 0 3236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5425
timestamp 1711653199
transform 1 0 3164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5426
timestamp 1711653199
transform 1 0 2876 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5427
timestamp 1711653199
transform 1 0 3316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5428
timestamp 1711653199
transform 1 0 3252 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5429
timestamp 1711653199
transform 1 0 3268 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5430
timestamp 1711653199
transform 1 0 3188 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5431
timestamp 1711653199
transform 1 0 3396 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_5432
timestamp 1711653199
transform 1 0 3396 0 1 1645
box -2 -2 2 2
use M2_M1  M2_M1_5433
timestamp 1711653199
transform 1 0 3372 0 1 1645
box -2 -2 2 2
use M2_M1  M2_M1_5434
timestamp 1711653199
transform 1 0 3372 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5435
timestamp 1711653199
transform 1 0 3356 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5436
timestamp 1711653199
transform 1 0 3132 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5437
timestamp 1711653199
transform 1 0 3396 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5438
timestamp 1711653199
transform 1 0 3348 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5439
timestamp 1711653199
transform 1 0 2820 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5440
timestamp 1711653199
transform 1 0 2724 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5441
timestamp 1711653199
transform 1 0 2700 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5442
timestamp 1711653199
transform 1 0 2508 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5443
timestamp 1711653199
transform 1 0 3132 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5444
timestamp 1711653199
transform 1 0 2844 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5445
timestamp 1711653199
transform 1 0 2772 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5446
timestamp 1711653199
transform 1 0 2436 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_5447
timestamp 1711653199
transform 1 0 2764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_5448
timestamp 1711653199
transform 1 0 2708 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5449
timestamp 1711653199
transform 1 0 2692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5450
timestamp 1711653199
transform 1 0 2684 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_5451
timestamp 1711653199
transform 1 0 2700 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_5452
timestamp 1711653199
transform 1 0 2628 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_5453
timestamp 1711653199
transform 1 0 2868 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5454
timestamp 1711653199
transform 1 0 2852 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_5455
timestamp 1711653199
transform 1 0 2844 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5456
timestamp 1711653199
transform 1 0 2780 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5457
timestamp 1711653199
transform 1 0 2764 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_5458
timestamp 1711653199
transform 1 0 2908 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5459
timestamp 1711653199
transform 1 0 2860 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_5460
timestamp 1711653199
transform 1 0 2756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5461
timestamp 1711653199
transform 1 0 2636 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5462
timestamp 1711653199
transform 1 0 2764 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5463
timestamp 1711653199
transform 1 0 2756 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5464
timestamp 1711653199
transform 1 0 2748 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5465
timestamp 1711653199
transform 1 0 2740 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5466
timestamp 1711653199
transform 1 0 2620 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_5467
timestamp 1711653199
transform 1 0 2716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_5468
timestamp 1711653199
transform 1 0 2708 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_5469
timestamp 1711653199
transform 1 0 2708 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5470
timestamp 1711653199
transform 1 0 2700 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_5471
timestamp 1711653199
transform 1 0 2980 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_5472
timestamp 1711653199
transform 1 0 2940 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5473
timestamp 1711653199
transform 1 0 2924 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5474
timestamp 1711653199
transform 1 0 2916 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_5475
timestamp 1711653199
transform 1 0 2860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5476
timestamp 1711653199
transform 1 0 2724 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_5477
timestamp 1711653199
transform 1 0 2724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5478
timestamp 1711653199
transform 1 0 3028 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5479
timestamp 1711653199
transform 1 0 3028 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5480
timestamp 1711653199
transform 1 0 3004 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5481
timestamp 1711653199
transform 1 0 2892 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5482
timestamp 1711653199
transform 1 0 2788 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5483
timestamp 1711653199
transform 1 0 2644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5484
timestamp 1711653199
transform 1 0 2636 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_5485
timestamp 1711653199
transform 1 0 2468 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5486
timestamp 1711653199
transform 1 0 2820 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5487
timestamp 1711653199
transform 1 0 2748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_5488
timestamp 1711653199
transform 1 0 3156 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5489
timestamp 1711653199
transform 1 0 2988 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5490
timestamp 1711653199
transform 1 0 2988 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_5491
timestamp 1711653199
transform 1 0 3148 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5492
timestamp 1711653199
transform 1 0 3004 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5493
timestamp 1711653199
transform 1 0 2852 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_5494
timestamp 1711653199
transform 1 0 2780 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_5495
timestamp 1711653199
transform 1 0 2748 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_5496
timestamp 1711653199
transform 1 0 2732 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_5497
timestamp 1711653199
transform 1 0 2876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5498
timestamp 1711653199
transform 1 0 2692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_5499
timestamp 1711653199
transform 1 0 3228 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5500
timestamp 1711653199
transform 1 0 2916 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5501
timestamp 1711653199
transform 1 0 2916 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5502
timestamp 1711653199
transform 1 0 2916 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5503
timestamp 1711653199
transform 1 0 2844 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5504
timestamp 1711653199
transform 1 0 2732 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5505
timestamp 1711653199
transform 1 0 2732 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5506
timestamp 1711653199
transform 1 0 2780 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_5507
timestamp 1711653199
transform 1 0 2740 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_5508
timestamp 1711653199
transform 1 0 2804 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5509
timestamp 1711653199
transform 1 0 2740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5510
timestamp 1711653199
transform 1 0 2708 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5511
timestamp 1711653199
transform 1 0 2436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5512
timestamp 1711653199
transform 1 0 2956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5513
timestamp 1711653199
transform 1 0 2892 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5514
timestamp 1711653199
transform 1 0 2556 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5515
timestamp 1711653199
transform 1 0 2340 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5516
timestamp 1711653199
transform 1 0 2516 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5517
timestamp 1711653199
transform 1 0 2508 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5518
timestamp 1711653199
transform 1 0 2500 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5519
timestamp 1711653199
transform 1 0 2484 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5520
timestamp 1711653199
transform 1 0 2444 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5521
timestamp 1711653199
transform 1 0 2412 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5522
timestamp 1711653199
transform 1 0 2812 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5523
timestamp 1711653199
transform 1 0 2772 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5524
timestamp 1711653199
transform 1 0 2812 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5525
timestamp 1711653199
transform 1 0 2748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5526
timestamp 1711653199
transform 1 0 2748 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5527
timestamp 1711653199
transform 1 0 2348 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5528
timestamp 1711653199
transform 1 0 2716 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5529
timestamp 1711653199
transform 1 0 2700 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5530
timestamp 1711653199
transform 1 0 2772 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5531
timestamp 1711653199
transform 1 0 2732 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5532
timestamp 1711653199
transform 1 0 2740 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5533
timestamp 1711653199
transform 1 0 2732 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5534
timestamp 1711653199
transform 1 0 2780 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5535
timestamp 1711653199
transform 1 0 2748 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5536
timestamp 1711653199
transform 1 0 2772 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5537
timestamp 1711653199
transform 1 0 2700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5538
timestamp 1711653199
transform 1 0 2724 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5539
timestamp 1711653199
transform 1 0 2668 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5540
timestamp 1711653199
transform 1 0 2628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5541
timestamp 1711653199
transform 1 0 2516 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5542
timestamp 1711653199
transform 1 0 2740 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5543
timestamp 1711653199
transform 1 0 2716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5544
timestamp 1711653199
transform 1 0 2716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5545
timestamp 1711653199
transform 1 0 2692 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5546
timestamp 1711653199
transform 1 0 2668 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5547
timestamp 1711653199
transform 1 0 2612 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5548
timestamp 1711653199
transform 1 0 2812 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5549
timestamp 1711653199
transform 1 0 2804 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5550
timestamp 1711653199
transform 1 0 2732 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_5551
timestamp 1711653199
transform 1 0 2596 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5552
timestamp 1711653199
transform 1 0 2692 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5553
timestamp 1711653199
transform 1 0 2684 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5554
timestamp 1711653199
transform 1 0 2700 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5555
timestamp 1711653199
transform 1 0 2564 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5556
timestamp 1711653199
transform 1 0 2244 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5557
timestamp 1711653199
transform 1 0 2236 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5558
timestamp 1711653199
transform 1 0 2692 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5559
timestamp 1711653199
transform 1 0 2636 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5560
timestamp 1711653199
transform 1 0 2652 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5561
timestamp 1711653199
transform 1 0 2652 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5562
timestamp 1711653199
transform 1 0 2460 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5563
timestamp 1711653199
transform 1 0 2356 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5564
timestamp 1711653199
transform 1 0 3012 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5565
timestamp 1711653199
transform 1 0 2820 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_5566
timestamp 1711653199
transform 1 0 2652 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5567
timestamp 1711653199
transform 1 0 2636 0 1 1734
box -2 -2 2 2
use M2_M1  M2_M1_5568
timestamp 1711653199
transform 1 0 2700 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5569
timestamp 1711653199
transform 1 0 2620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5570
timestamp 1711653199
transform 1 0 2604 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5571
timestamp 1711653199
transform 1 0 2604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5572
timestamp 1711653199
transform 1 0 2844 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5573
timestamp 1711653199
transform 1 0 2844 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5574
timestamp 1711653199
transform 1 0 2812 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5575
timestamp 1711653199
transform 1 0 2636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5576
timestamp 1711653199
transform 1 0 2636 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5577
timestamp 1711653199
transform 1 0 2644 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5578
timestamp 1711653199
transform 1 0 2572 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5579
timestamp 1711653199
transform 1 0 2588 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5580
timestamp 1711653199
transform 1 0 2356 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5581
timestamp 1711653199
transform 1 0 2652 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5582
timestamp 1711653199
transform 1 0 2636 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_5583
timestamp 1711653199
transform 1 0 2500 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5584
timestamp 1711653199
transform 1 0 2492 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5585
timestamp 1711653199
transform 1 0 2468 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5586
timestamp 1711653199
transform 1 0 2396 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5587
timestamp 1711653199
transform 1 0 2660 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5588
timestamp 1711653199
transform 1 0 2452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5589
timestamp 1711653199
transform 1 0 2940 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5590
timestamp 1711653199
transform 1 0 2460 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5591
timestamp 1711653199
transform 1 0 2940 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5592
timestamp 1711653199
transform 1 0 2900 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5593
timestamp 1711653199
transform 1 0 2812 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_5594
timestamp 1711653199
transform 1 0 2716 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5595
timestamp 1711653199
transform 1 0 2940 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5596
timestamp 1711653199
transform 1 0 2844 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5597
timestamp 1711653199
transform 1 0 2932 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5598
timestamp 1711653199
transform 1 0 2828 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5599
timestamp 1711653199
transform 1 0 3004 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5600
timestamp 1711653199
transform 1 0 2996 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5601
timestamp 1711653199
transform 1 0 2956 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_5602
timestamp 1711653199
transform 1 0 2868 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5603
timestamp 1711653199
transform 1 0 2812 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5604
timestamp 1711653199
transform 1 0 3108 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5605
timestamp 1711653199
transform 1 0 2972 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5606
timestamp 1711653199
transform 1 0 2932 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_5607
timestamp 1711653199
transform 1 0 2900 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5608
timestamp 1711653199
transform 1 0 2884 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_5609
timestamp 1711653199
transform 1 0 2884 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5610
timestamp 1711653199
transform 1 0 2700 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5611
timestamp 1711653199
transform 1 0 2660 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_5612
timestamp 1711653199
transform 1 0 2660 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_5613
timestamp 1711653199
transform 1 0 2660 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5614
timestamp 1711653199
transform 1 0 2644 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5615
timestamp 1711653199
transform 1 0 2644 0 1 1585
box -2 -2 2 2
use M2_M1  M2_M1_5616
timestamp 1711653199
transform 1 0 2692 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_5617
timestamp 1711653199
transform 1 0 2564 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5618
timestamp 1711653199
transform 1 0 2604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5619
timestamp 1711653199
transform 1 0 2532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5620
timestamp 1711653199
transform 1 0 2572 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5621
timestamp 1711653199
transform 1 0 2516 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5622
timestamp 1711653199
transform 1 0 2508 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5623
timestamp 1711653199
transform 1 0 2644 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5624
timestamp 1711653199
transform 1 0 2572 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5625
timestamp 1711653199
transform 1 0 2596 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5626
timestamp 1711653199
transform 1 0 2524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5627
timestamp 1711653199
transform 1 0 2644 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5628
timestamp 1711653199
transform 1 0 2556 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5629
timestamp 1711653199
transform 1 0 2668 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5630
timestamp 1711653199
transform 1 0 2668 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5631
timestamp 1711653199
transform 1 0 2580 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5632
timestamp 1711653199
transform 1 0 2444 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5633
timestamp 1711653199
transform 1 0 2660 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5634
timestamp 1711653199
transform 1 0 2580 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5635
timestamp 1711653199
transform 1 0 2564 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5636
timestamp 1711653199
transform 1 0 2564 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5637
timestamp 1711653199
transform 1 0 2660 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5638
timestamp 1711653199
transform 1 0 2540 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5639
timestamp 1711653199
transform 1 0 2556 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5640
timestamp 1711653199
transform 1 0 2460 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5641
timestamp 1711653199
transform 1 0 2668 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5642
timestamp 1711653199
transform 1 0 2652 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5643
timestamp 1711653199
transform 1 0 2916 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5644
timestamp 1711653199
transform 1 0 2484 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5645
timestamp 1711653199
transform 1 0 2892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5646
timestamp 1711653199
transform 1 0 2892 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5647
timestamp 1711653199
transform 1 0 2940 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5648
timestamp 1711653199
transform 1 0 2892 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5649
timestamp 1711653199
transform 1 0 2916 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5650
timestamp 1711653199
transform 1 0 2852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5651
timestamp 1711653199
transform 1 0 2900 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_5652
timestamp 1711653199
transform 1 0 2892 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5653
timestamp 1711653199
transform 1 0 2828 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_5654
timestamp 1711653199
transform 1 0 2796 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5655
timestamp 1711653199
transform 1 0 2772 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5656
timestamp 1711653199
transform 1 0 2756 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5657
timestamp 1711653199
transform 1 0 2788 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5658
timestamp 1711653199
transform 1 0 2788 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5659
timestamp 1711653199
transform 1 0 2732 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5660
timestamp 1711653199
transform 1 0 2724 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5661
timestamp 1711653199
transform 1 0 2940 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5662
timestamp 1711653199
transform 1 0 2724 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5663
timestamp 1711653199
transform 1 0 2756 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5664
timestamp 1711653199
transform 1 0 2452 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5665
timestamp 1711653199
transform 1 0 2516 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5666
timestamp 1711653199
transform 1 0 2484 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5667
timestamp 1711653199
transform 1 0 2940 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5668
timestamp 1711653199
transform 1 0 2860 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5669
timestamp 1711653199
transform 1 0 2876 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5670
timestamp 1711653199
transform 1 0 2868 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5671
timestamp 1711653199
transform 1 0 2764 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5672
timestamp 1711653199
transform 1 0 2396 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5673
timestamp 1711653199
transform 1 0 2852 0 1 1685
box -2 -2 2 2
use M2_M1  M2_M1_5674
timestamp 1711653199
transform 1 0 2852 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5675
timestamp 1711653199
transform 1 0 2820 0 1 1685
box -2 -2 2 2
use M2_M1  M2_M1_5676
timestamp 1711653199
transform 1 0 2796 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5677
timestamp 1711653199
transform 1 0 2764 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5678
timestamp 1711653199
transform 1 0 2764 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5679
timestamp 1711653199
transform 1 0 2940 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5680
timestamp 1711653199
transform 1 0 2740 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5681
timestamp 1711653199
transform 1 0 2700 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5682
timestamp 1711653199
transform 1 0 2420 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5683
timestamp 1711653199
transform 1 0 2916 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5684
timestamp 1711653199
transform 1 0 2916 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5685
timestamp 1711653199
transform 1 0 3316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5686
timestamp 1711653199
transform 1 0 3140 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5687
timestamp 1711653199
transform 1 0 3132 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5688
timestamp 1711653199
transform 1 0 3084 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5689
timestamp 1711653199
transform 1 0 3036 0 1 1555
box -2 -2 2 2
use M2_M1  M2_M1_5690
timestamp 1711653199
transform 1 0 2996 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5691
timestamp 1711653199
transform 1 0 3116 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_5692
timestamp 1711653199
transform 1 0 2436 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5693
timestamp 1711653199
transform 1 0 3108 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5694
timestamp 1711653199
transform 1 0 3076 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5695
timestamp 1711653199
transform 1 0 3076 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5696
timestamp 1711653199
transform 1 0 3036 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_5697
timestamp 1711653199
transform 1 0 3028 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_5698
timestamp 1711653199
transform 1 0 3028 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5699
timestamp 1711653199
transform 1 0 3012 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_5700
timestamp 1711653199
transform 1 0 3004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_5701
timestamp 1711653199
transform 1 0 3084 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_5702
timestamp 1711653199
transform 1 0 3012 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_5703
timestamp 1711653199
transform 1 0 3068 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_5704
timestamp 1711653199
transform 1 0 2948 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_5705
timestamp 1711653199
transform 1 0 3092 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5706
timestamp 1711653199
transform 1 0 3084 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5707
timestamp 1711653199
transform 1 0 3052 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5708
timestamp 1711653199
transform 1 0 3028 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_5709
timestamp 1711653199
transform 1 0 3068 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5710
timestamp 1711653199
transform 1 0 3068 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5711
timestamp 1711653199
transform 1 0 2940 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5712
timestamp 1711653199
transform 1 0 3084 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5713
timestamp 1711653199
transform 1 0 3084 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5714
timestamp 1711653199
transform 1 0 3084 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5715
timestamp 1711653199
transform 1 0 3060 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5716
timestamp 1711653199
transform 1 0 3108 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5717
timestamp 1711653199
transform 1 0 2972 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5718
timestamp 1711653199
transform 1 0 3052 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5719
timestamp 1711653199
transform 1 0 2956 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5720
timestamp 1711653199
transform 1 0 3020 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5721
timestamp 1711653199
transform 1 0 3020 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5722
timestamp 1711653199
transform 1 0 3012 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5723
timestamp 1711653199
transform 1 0 2956 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5724
timestamp 1711653199
transform 1 0 2820 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5725
timestamp 1711653199
transform 1 0 2964 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_5726
timestamp 1711653199
transform 1 0 2956 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5727
timestamp 1711653199
transform 1 0 3172 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5728
timestamp 1711653199
transform 1 0 3132 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5729
timestamp 1711653199
transform 1 0 3100 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5730
timestamp 1711653199
transform 1 0 3020 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5731
timestamp 1711653199
transform 1 0 2988 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_5732
timestamp 1711653199
transform 1 0 3132 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_5733
timestamp 1711653199
transform 1 0 3108 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5734
timestamp 1711653199
transform 1 0 3084 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5735
timestamp 1711653199
transform 1 0 3068 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5736
timestamp 1711653199
transform 1 0 3356 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5737
timestamp 1711653199
transform 1 0 3324 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5738
timestamp 1711653199
transform 1 0 3332 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5739
timestamp 1711653199
transform 1 0 3292 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5740
timestamp 1711653199
transform 1 0 3188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5741
timestamp 1711653199
transform 1 0 3364 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5742
timestamp 1711653199
transform 1 0 3356 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5743
timestamp 1711653199
transform 1 0 3332 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5744
timestamp 1711653199
transform 1 0 3332 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5745
timestamp 1711653199
transform 1 0 3348 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5746
timestamp 1711653199
transform 1 0 3348 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5747
timestamp 1711653199
transform 1 0 3332 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_5748
timestamp 1711653199
transform 1 0 3308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5749
timestamp 1711653199
transform 1 0 3276 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5750
timestamp 1711653199
transform 1 0 3380 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_5751
timestamp 1711653199
transform 1 0 3364 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5752
timestamp 1711653199
transform 1 0 3388 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_5753
timestamp 1711653199
transform 1 0 3356 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_5754
timestamp 1711653199
transform 1 0 3332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_5755
timestamp 1711653199
transform 1 0 2756 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_5756
timestamp 1711653199
transform 1 0 2732 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5757
timestamp 1711653199
transform 1 0 3260 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5758
timestamp 1711653199
transform 1 0 3156 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5759
timestamp 1711653199
transform 1 0 3076 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5760
timestamp 1711653199
transform 1 0 2892 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5761
timestamp 1711653199
transform 1 0 2748 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5762
timestamp 1711653199
transform 1 0 2748 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5763
timestamp 1711653199
transform 1 0 3284 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5764
timestamp 1711653199
transform 1 0 3172 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5765
timestamp 1711653199
transform 1 0 3108 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5766
timestamp 1711653199
transform 1 0 2908 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5767
timestamp 1711653199
transform 1 0 2780 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5768
timestamp 1711653199
transform 1 0 2780 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5769
timestamp 1711653199
transform 1 0 2764 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5770
timestamp 1711653199
transform 1 0 2764 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5771
timestamp 1711653199
transform 1 0 2932 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_5772
timestamp 1711653199
transform 1 0 2900 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5773
timestamp 1711653199
transform 1 0 3132 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5774
timestamp 1711653199
transform 1 0 3100 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5775
timestamp 1711653199
transform 1 0 3172 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_5776
timestamp 1711653199
transform 1 0 3164 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5777
timestamp 1711653199
transform 1 0 3292 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5778
timestamp 1711653199
transform 1 0 3284 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5779
timestamp 1711653199
transform 1 0 3276 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_5780
timestamp 1711653199
transform 1 0 3300 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5781
timestamp 1711653199
transform 1 0 3300 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5782
timestamp 1711653199
transform 1 0 3292 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_5783
timestamp 1711653199
transform 1 0 3332 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5784
timestamp 1711653199
transform 1 0 3300 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5785
timestamp 1711653199
transform 1 0 3324 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5786
timestamp 1711653199
transform 1 0 3244 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5787
timestamp 1711653199
transform 1 0 3244 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5788
timestamp 1711653199
transform 1 0 3340 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5789
timestamp 1711653199
transform 1 0 3324 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5790
timestamp 1711653199
transform 1 0 3300 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_5791
timestamp 1711653199
transform 1 0 3268 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5792
timestamp 1711653199
transform 1 0 3348 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_5793
timestamp 1711653199
transform 1 0 3180 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5794
timestamp 1711653199
transform 1 0 3340 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_5795
timestamp 1711653199
transform 1 0 3324 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_5796
timestamp 1711653199
transform 1 0 3340 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_5797
timestamp 1711653199
transform 1 0 3316 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5798
timestamp 1711653199
transform 1 0 3244 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_5799
timestamp 1711653199
transform 1 0 3236 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5800
timestamp 1711653199
transform 1 0 3260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5801
timestamp 1711653199
transform 1 0 3180 0 1 2305
box -2 -2 2 2
use M2_M1  M2_M1_5802
timestamp 1711653199
transform 1 0 3180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5803
timestamp 1711653199
transform 1 0 3252 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_5804
timestamp 1711653199
transform 1 0 3212 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5805
timestamp 1711653199
transform 1 0 3260 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5806
timestamp 1711653199
transform 1 0 3188 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5807
timestamp 1711653199
transform 1 0 3268 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5808
timestamp 1711653199
transform 1 0 3188 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5809
timestamp 1711653199
transform 1 0 3220 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5810
timestamp 1711653199
transform 1 0 3204 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5811
timestamp 1711653199
transform 1 0 2796 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5812
timestamp 1711653199
transform 1 0 2788 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5813
timestamp 1711653199
transform 1 0 2676 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_5814
timestamp 1711653199
transform 1 0 2020 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5815
timestamp 1711653199
transform 1 0 2020 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5816
timestamp 1711653199
transform 1 0 2436 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5817
timestamp 1711653199
transform 1 0 2420 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5818
timestamp 1711653199
transform 1 0 2316 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5819
timestamp 1711653199
transform 1 0 2212 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5820
timestamp 1711653199
transform 1 0 2148 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5821
timestamp 1711653199
transform 1 0 2124 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5822
timestamp 1711653199
transform 1 0 2300 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5823
timestamp 1711653199
transform 1 0 2300 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5824
timestamp 1711653199
transform 1 0 2740 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5825
timestamp 1711653199
transform 1 0 2636 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5826
timestamp 1711653199
transform 1 0 2532 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5827
timestamp 1711653199
transform 1 0 2492 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5828
timestamp 1711653199
transform 1 0 1964 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5829
timestamp 1711653199
transform 1 0 1948 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5830
timestamp 1711653199
transform 1 0 1908 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5831
timestamp 1711653199
transform 1 0 1860 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5832
timestamp 1711653199
transform 1 0 1660 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5833
timestamp 1711653199
transform 1 0 1620 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5834
timestamp 1711653199
transform 1 0 1756 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5835
timestamp 1711653199
transform 1 0 1740 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5836
timestamp 1711653199
transform 1 0 1492 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5837
timestamp 1711653199
transform 1 0 1492 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5838
timestamp 1711653199
transform 1 0 1324 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5839
timestamp 1711653199
transform 1 0 1284 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5840
timestamp 1711653199
transform 1 0 964 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5841
timestamp 1711653199
transform 1 0 868 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5842
timestamp 1711653199
transform 1 0 788 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5843
timestamp 1711653199
transform 1 0 628 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5844
timestamp 1711653199
transform 1 0 1108 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5845
timestamp 1711653199
transform 1 0 1044 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5846
timestamp 1711653199
transform 1 0 748 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5847
timestamp 1711653199
transform 1 0 740 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5848
timestamp 1711653199
transform 1 0 452 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5849
timestamp 1711653199
transform 1 0 404 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5850
timestamp 1711653199
transform 1 0 404 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5851
timestamp 1711653199
transform 1 0 308 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5852
timestamp 1711653199
transform 1 0 300 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5853
timestamp 1711653199
transform 1 0 284 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5854
timestamp 1711653199
transform 1 0 220 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5855
timestamp 1711653199
transform 1 0 140 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5856
timestamp 1711653199
transform 1 0 220 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5857
timestamp 1711653199
transform 1 0 132 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_5858
timestamp 1711653199
transform 1 0 180 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5859
timestamp 1711653199
transform 1 0 132 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_5860
timestamp 1711653199
transform 1 0 228 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5861
timestamp 1711653199
transform 1 0 204 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5862
timestamp 1711653199
transform 1 0 508 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5863
timestamp 1711653199
transform 1 0 468 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_5864
timestamp 1711653199
transform 1 0 372 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5865
timestamp 1711653199
transform 1 0 372 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5866
timestamp 1711653199
transform 1 0 756 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5867
timestamp 1711653199
transform 1 0 716 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5868
timestamp 1711653199
transform 1 0 1004 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5869
timestamp 1711653199
transform 1 0 964 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_5870
timestamp 1711653199
transform 1 0 1532 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5871
timestamp 1711653199
transform 1 0 1524 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5872
timestamp 1711653199
transform 1 0 1804 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5873
timestamp 1711653199
transform 1 0 1804 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_5874
timestamp 1711653199
transform 1 0 1884 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_5875
timestamp 1711653199
transform 1 0 1844 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_5876
timestamp 1711653199
transform 1 0 2012 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_5877
timestamp 1711653199
transform 1 0 2004 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_5878
timestamp 1711653199
transform 1 0 2828 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5879
timestamp 1711653199
transform 1 0 2804 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5880
timestamp 1711653199
transform 1 0 2652 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5881
timestamp 1711653199
transform 1 0 2628 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_5882
timestamp 1711653199
transform 1 0 2660 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5883
timestamp 1711653199
transform 1 0 2644 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5884
timestamp 1711653199
transform 1 0 2636 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_5885
timestamp 1711653199
transform 1 0 2580 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5886
timestamp 1711653199
transform 1 0 2532 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_5887
timestamp 1711653199
transform 1 0 2684 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5888
timestamp 1711653199
transform 1 0 2652 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_5889
timestamp 1711653199
transform 1 0 2748 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5890
timestamp 1711653199
transform 1 0 2628 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5891
timestamp 1711653199
transform 1 0 2556 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5892
timestamp 1711653199
transform 1 0 2668 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5893
timestamp 1711653199
transform 1 0 2652 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_5894
timestamp 1711653199
transform 1 0 2668 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5895
timestamp 1711653199
transform 1 0 2652 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5896
timestamp 1711653199
transform 1 0 2116 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5897
timestamp 1711653199
transform 1 0 2100 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_5898
timestamp 1711653199
transform 1 0 2540 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5899
timestamp 1711653199
transform 1 0 2484 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5900
timestamp 1711653199
transform 1 0 2404 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5901
timestamp 1711653199
transform 1 0 2380 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5902
timestamp 1711653199
transform 1 0 2404 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5903
timestamp 1711653199
transform 1 0 2372 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5904
timestamp 1711653199
transform 1 0 2364 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5905
timestamp 1711653199
transform 1 0 2340 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5906
timestamp 1711653199
transform 1 0 2540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5907
timestamp 1711653199
transform 1 0 2508 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5908
timestamp 1711653199
transform 1 0 2476 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5909
timestamp 1711653199
transform 1 0 2468 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5910
timestamp 1711653199
transform 1 0 2196 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5911
timestamp 1711653199
transform 1 0 2196 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5912
timestamp 1711653199
transform 1 0 2516 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5913
timestamp 1711653199
transform 1 0 2268 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5914
timestamp 1711653199
transform 1 0 2244 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5915
timestamp 1711653199
transform 1 0 2108 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5916
timestamp 1711653199
transform 1 0 2084 0 1 2985
box -2 -2 2 2
use M2_M1  M2_M1_5917
timestamp 1711653199
transform 1 0 2012 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5918
timestamp 1711653199
transform 1 0 1684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5919
timestamp 1711653199
transform 1 0 2420 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5920
timestamp 1711653199
transform 1 0 2244 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5921
timestamp 1711653199
transform 1 0 2612 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5922
timestamp 1711653199
transform 1 0 2444 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5923
timestamp 1711653199
transform 1 0 2396 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5924
timestamp 1711653199
transform 1 0 2484 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5925
timestamp 1711653199
transform 1 0 2452 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_5926
timestamp 1711653199
transform 1 0 2468 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5927
timestamp 1711653199
transform 1 0 2348 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5928
timestamp 1711653199
transform 1 0 2228 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5929
timestamp 1711653199
transform 1 0 2204 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5930
timestamp 1711653199
transform 1 0 1516 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5931
timestamp 1711653199
transform 1 0 1516 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5932
timestamp 1711653199
transform 1 0 2284 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5933
timestamp 1711653199
transform 1 0 2180 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5934
timestamp 1711653199
transform 1 0 1380 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5935
timestamp 1711653199
transform 1 0 2388 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5936
timestamp 1711653199
transform 1 0 2316 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5937
timestamp 1711653199
transform 1 0 2396 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_5938
timestamp 1711653199
transform 1 0 2364 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5939
timestamp 1711653199
transform 1 0 2340 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5940
timestamp 1711653199
transform 1 0 2340 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5941
timestamp 1711653199
transform 1 0 2252 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_5942
timestamp 1711653199
transform 1 0 2124 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5943
timestamp 1711653199
transform 1 0 1980 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5944
timestamp 1711653199
transform 1 0 2276 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_5945
timestamp 1711653199
transform 1 0 2260 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5946
timestamp 1711653199
transform 1 0 3132 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5947
timestamp 1711653199
transform 1 0 2732 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_5948
timestamp 1711653199
transform 1 0 2644 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5949
timestamp 1711653199
transform 1 0 1420 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5950
timestamp 1711653199
transform 1 0 1372 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_5951
timestamp 1711653199
transform 1 0 1388 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5952
timestamp 1711653199
transform 1 0 1180 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5953
timestamp 1711653199
transform 1 0 1124 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5954
timestamp 1711653199
transform 1 0 1124 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5955
timestamp 1711653199
transform 1 0 1124 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_5956
timestamp 1711653199
transform 1 0 1100 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5957
timestamp 1711653199
transform 1 0 1044 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5958
timestamp 1711653199
transform 1 0 1196 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5959
timestamp 1711653199
transform 1 0 1172 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5960
timestamp 1711653199
transform 1 0 1132 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5961
timestamp 1711653199
transform 1 0 1108 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_5962
timestamp 1711653199
transform 1 0 972 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5963
timestamp 1711653199
transform 1 0 916 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5964
timestamp 1711653199
transform 1 0 844 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_5965
timestamp 1711653199
transform 1 0 1268 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_5966
timestamp 1711653199
transform 1 0 1268 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_5967
timestamp 1711653199
transform 1 0 1252 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_5968
timestamp 1711653199
transform 1 0 1212 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_5969
timestamp 1711653199
transform 1 0 1196 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_5970
timestamp 1711653199
transform 1 0 1188 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_5971
timestamp 1711653199
transform 1 0 1172 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_5972
timestamp 1711653199
transform 1 0 1396 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5973
timestamp 1711653199
transform 1 0 1316 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5974
timestamp 1711653199
transform 1 0 1252 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5975
timestamp 1711653199
transform 1 0 1164 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5976
timestamp 1711653199
transform 1 0 1492 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5977
timestamp 1711653199
transform 1 0 1404 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5978
timestamp 1711653199
transform 1 0 1324 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5979
timestamp 1711653199
transform 1 0 1188 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5980
timestamp 1711653199
transform 1 0 900 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5981
timestamp 1711653199
transform 1 0 780 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5982
timestamp 1711653199
transform 1 0 756 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5983
timestamp 1711653199
transform 1 0 1460 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_5984
timestamp 1711653199
transform 1 0 1428 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5985
timestamp 1711653199
transform 1 0 2044 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_5986
timestamp 1711653199
transform 1 0 2012 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5987
timestamp 1711653199
transform 1 0 1660 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5988
timestamp 1711653199
transform 1 0 1524 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_5989
timestamp 1711653199
transform 1 0 1364 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_5990
timestamp 1711653199
transform 1 0 1844 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_5991
timestamp 1711653199
transform 1 0 1820 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5992
timestamp 1711653199
transform 1 0 1764 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_5993
timestamp 1711653199
transform 1 0 1748 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5994
timestamp 1711653199
transform 1 0 1884 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_5995
timestamp 1711653199
transform 1 0 1796 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_5996
timestamp 1711653199
transform 1 0 1732 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_5997
timestamp 1711653199
transform 1 0 1668 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_5998
timestamp 1711653199
transform 1 0 1588 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_5999
timestamp 1711653199
transform 1 0 1540 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6000
timestamp 1711653199
transform 1 0 1460 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6001
timestamp 1711653199
transform 1 0 1332 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6002
timestamp 1711653199
transform 1 0 1652 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6003
timestamp 1711653199
transform 1 0 1612 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6004
timestamp 1711653199
transform 1 0 1780 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6005
timestamp 1711653199
transform 1 0 1636 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6006
timestamp 1711653199
transform 1 0 1732 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6007
timestamp 1711653199
transform 1 0 1724 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6008
timestamp 1711653199
transform 1 0 1844 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6009
timestamp 1711653199
transform 1 0 1708 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6010
timestamp 1711653199
transform 1 0 1572 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6011
timestamp 1711653199
transform 1 0 1492 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6012
timestamp 1711653199
transform 1 0 1524 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6013
timestamp 1711653199
transform 1 0 1492 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6014
timestamp 1711653199
transform 1 0 1564 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6015
timestamp 1711653199
transform 1 0 1548 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6016
timestamp 1711653199
transform 1 0 1524 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6017
timestamp 1711653199
transform 1 0 1436 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6018
timestamp 1711653199
transform 1 0 1396 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6019
timestamp 1711653199
transform 1 0 1380 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6020
timestamp 1711653199
transform 1 0 1364 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6021
timestamp 1711653199
transform 1 0 1340 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6022
timestamp 1711653199
transform 1 0 1228 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6023
timestamp 1711653199
transform 1 0 1972 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6024
timestamp 1711653199
transform 1 0 1484 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6025
timestamp 1711653199
transform 1 0 1444 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6026
timestamp 1711653199
transform 1 0 1412 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6027
timestamp 1711653199
transform 1 0 1308 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6028
timestamp 1711653199
transform 1 0 1428 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6029
timestamp 1711653199
transform 1 0 1420 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6030
timestamp 1711653199
transform 1 0 1388 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6031
timestamp 1711653199
transform 1 0 1252 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6032
timestamp 1711653199
transform 1 0 1244 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6033
timestamp 1711653199
transform 1 0 1100 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6034
timestamp 1711653199
transform 1 0 1508 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6035
timestamp 1711653199
transform 1 0 1396 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6036
timestamp 1711653199
transform 1 0 1396 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6037
timestamp 1711653199
transform 1 0 1268 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6038
timestamp 1711653199
transform 1 0 1164 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6039
timestamp 1711653199
transform 1 0 1036 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6040
timestamp 1711653199
transform 1 0 964 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6041
timestamp 1711653199
transform 1 0 1372 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6042
timestamp 1711653199
transform 1 0 1340 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6043
timestamp 1711653199
transform 1 0 1412 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6044
timestamp 1711653199
transform 1 0 1348 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6045
timestamp 1711653199
transform 1 0 1332 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6046
timestamp 1711653199
transform 1 0 1308 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6047
timestamp 1711653199
transform 1 0 1356 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6048
timestamp 1711653199
transform 1 0 1324 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6049
timestamp 1711653199
transform 1 0 1228 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6050
timestamp 1711653199
transform 1 0 1084 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6051
timestamp 1711653199
transform 1 0 996 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6052
timestamp 1711653199
transform 1 0 996 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6053
timestamp 1711653199
transform 1 0 1100 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6054
timestamp 1711653199
transform 1 0 1068 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6055
timestamp 1711653199
transform 1 0 1252 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6056
timestamp 1711653199
transform 1 0 1076 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6057
timestamp 1711653199
transform 1 0 1068 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6058
timestamp 1711653199
transform 1 0 1068 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6059
timestamp 1711653199
transform 1 0 1004 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6060
timestamp 1711653199
transform 1 0 948 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6061
timestamp 1711653199
transform 1 0 1236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6062
timestamp 1711653199
transform 1 0 980 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6063
timestamp 1711653199
transform 1 0 980 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6064
timestamp 1711653199
transform 1 0 980 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6065
timestamp 1711653199
transform 1 0 1220 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6066
timestamp 1711653199
transform 1 0 1188 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6067
timestamp 1711653199
transform 1 0 1380 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6068
timestamp 1711653199
transform 1 0 1196 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6069
timestamp 1711653199
transform 1 0 1212 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6070
timestamp 1711653199
transform 1 0 1204 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6071
timestamp 1711653199
transform 1 0 1180 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6072
timestamp 1711653199
transform 1 0 1140 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6073
timestamp 1711653199
transform 1 0 1108 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6074
timestamp 1711653199
transform 1 0 1012 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6075
timestamp 1711653199
transform 1 0 1036 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6076
timestamp 1711653199
transform 1 0 892 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6077
timestamp 1711653199
transform 1 0 868 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6078
timestamp 1711653199
transform 1 0 804 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6079
timestamp 1711653199
transform 1 0 748 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6080
timestamp 1711653199
transform 1 0 708 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6081
timestamp 1711653199
transform 1 0 1100 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6082
timestamp 1711653199
transform 1 0 836 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6083
timestamp 1711653199
transform 1 0 828 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6084
timestamp 1711653199
transform 1 0 764 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6085
timestamp 1711653199
transform 1 0 732 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6086
timestamp 1711653199
transform 1 0 692 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6087
timestamp 1711653199
transform 1 0 1028 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6088
timestamp 1711653199
transform 1 0 1004 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6089
timestamp 1711653199
transform 1 0 996 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6090
timestamp 1711653199
transform 1 0 724 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_6091
timestamp 1711653199
transform 1 0 604 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6092
timestamp 1711653199
transform 1 0 660 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6093
timestamp 1711653199
transform 1 0 628 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6094
timestamp 1711653199
transform 1 0 1020 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6095
timestamp 1711653199
transform 1 0 836 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6096
timestamp 1711653199
transform 1 0 628 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6097
timestamp 1711653199
transform 1 0 564 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6098
timestamp 1711653199
transform 1 0 540 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6099
timestamp 1711653199
transform 1 0 532 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6100
timestamp 1711653199
transform 1 0 860 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6101
timestamp 1711653199
transform 1 0 676 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6102
timestamp 1711653199
transform 1 0 580 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6103
timestamp 1711653199
transform 1 0 564 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6104
timestamp 1711653199
transform 1 0 796 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6105
timestamp 1711653199
transform 1 0 596 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6106
timestamp 1711653199
transform 1 0 452 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6107
timestamp 1711653199
transform 1 0 380 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6108
timestamp 1711653199
transform 1 0 556 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6109
timestamp 1711653199
transform 1 0 476 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6110
timestamp 1711653199
transform 1 0 700 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6111
timestamp 1711653199
transform 1 0 556 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6112
timestamp 1711653199
transform 1 0 404 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6113
timestamp 1711653199
transform 1 0 300 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6114
timestamp 1711653199
transform 1 0 588 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6115
timestamp 1711653199
transform 1 0 444 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6116
timestamp 1711653199
transform 1 0 740 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6117
timestamp 1711653199
transform 1 0 612 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6118
timestamp 1711653199
transform 1 0 948 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6119
timestamp 1711653199
transform 1 0 868 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6120
timestamp 1711653199
transform 1 0 844 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6121
timestamp 1711653199
transform 1 0 804 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6122
timestamp 1711653199
transform 1 0 940 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6123
timestamp 1711653199
transform 1 0 892 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6124
timestamp 1711653199
transform 1 0 636 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6125
timestamp 1711653199
transform 1 0 564 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6126
timestamp 1711653199
transform 1 0 516 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6127
timestamp 1711653199
transform 1 0 500 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6128
timestamp 1711653199
transform 1 0 980 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6129
timestamp 1711653199
transform 1 0 836 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6130
timestamp 1711653199
transform 1 0 716 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6131
timestamp 1711653199
transform 1 0 660 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6132
timestamp 1711653199
transform 1 0 636 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6133
timestamp 1711653199
transform 1 0 620 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6134
timestamp 1711653199
transform 1 0 628 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6135
timestamp 1711653199
transform 1 0 236 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_6136
timestamp 1711653199
transform 1 0 628 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6137
timestamp 1711653199
transform 1 0 604 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6138
timestamp 1711653199
transform 1 0 676 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6139
timestamp 1711653199
transform 1 0 612 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6140
timestamp 1711653199
transform 1 0 860 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6141
timestamp 1711653199
transform 1 0 844 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6142
timestamp 1711653199
transform 1 0 756 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6143
timestamp 1711653199
transform 1 0 692 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6144
timestamp 1711653199
transform 1 0 692 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6145
timestamp 1711653199
transform 1 0 652 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6146
timestamp 1711653199
transform 1 0 556 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6147
timestamp 1711653199
transform 1 0 436 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_6148
timestamp 1711653199
transform 1 0 556 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6149
timestamp 1711653199
transform 1 0 532 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6150
timestamp 1711653199
transform 1 0 636 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6151
timestamp 1711653199
transform 1 0 540 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6152
timestamp 1711653199
transform 1 0 476 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6153
timestamp 1711653199
transform 1 0 244 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_6154
timestamp 1711653199
transform 1 0 476 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6155
timestamp 1711653199
transform 1 0 436 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6156
timestamp 1711653199
transform 1 0 676 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6157
timestamp 1711653199
transform 1 0 452 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6158
timestamp 1711653199
transform 1 0 508 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6159
timestamp 1711653199
transform 1 0 260 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6160
timestamp 1711653199
transform 1 0 508 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6161
timestamp 1711653199
transform 1 0 484 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6162
timestamp 1711653199
transform 1 0 740 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6163
timestamp 1711653199
transform 1 0 492 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6164
timestamp 1711653199
transform 1 0 1060 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6165
timestamp 1711653199
transform 1 0 1028 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6166
timestamp 1711653199
transform 1 0 980 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6167
timestamp 1711653199
transform 1 0 948 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6168
timestamp 1711653199
transform 1 0 852 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6169
timestamp 1711653199
transform 1 0 828 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6170
timestamp 1711653199
transform 1 0 1092 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6171
timestamp 1711653199
transform 1 0 940 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6172
timestamp 1711653199
transform 1 0 900 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6173
timestamp 1711653199
transform 1 0 1188 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_6174
timestamp 1711653199
transform 1 0 988 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6175
timestamp 1711653199
transform 1 0 892 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_6176
timestamp 1711653199
transform 1 0 588 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6177
timestamp 1711653199
transform 1 0 564 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6178
timestamp 1711653199
transform 1 0 700 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6179
timestamp 1711653199
transform 1 0 628 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6180
timestamp 1711653199
transform 1 0 1020 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6181
timestamp 1711653199
transform 1 0 716 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6182
timestamp 1711653199
transform 1 0 1220 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_6183
timestamp 1711653199
transform 1 0 1012 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6184
timestamp 1711653199
transform 1 0 932 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6185
timestamp 1711653199
transform 1 0 844 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6186
timestamp 1711653199
transform 1 0 836 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6187
timestamp 1711653199
transform 1 0 796 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6188
timestamp 1711653199
transform 1 0 572 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6189
timestamp 1711653199
transform 1 0 404 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6190
timestamp 1711653199
transform 1 0 668 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6191
timestamp 1711653199
transform 1 0 604 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6192
timestamp 1711653199
transform 1 0 804 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6193
timestamp 1711653199
transform 1 0 668 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6194
timestamp 1711653199
transform 1 0 748 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6195
timestamp 1711653199
transform 1 0 740 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6196
timestamp 1711653199
transform 1 0 844 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6197
timestamp 1711653199
transform 1 0 748 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6198
timestamp 1711653199
transform 1 0 956 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6199
timestamp 1711653199
transform 1 0 916 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6200
timestamp 1711653199
transform 1 0 940 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6201
timestamp 1711653199
transform 1 0 916 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6202
timestamp 1711653199
transform 1 0 1316 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6203
timestamp 1711653199
transform 1 0 1252 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6204
timestamp 1711653199
transform 1 0 1196 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6205
timestamp 1711653199
transform 1 0 1084 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6206
timestamp 1711653199
transform 1 0 1060 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_6207
timestamp 1711653199
transform 1 0 1052 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6208
timestamp 1711653199
transform 1 0 1292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6209
timestamp 1711653199
transform 1 0 1284 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6210
timestamp 1711653199
transform 1 0 1220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6211
timestamp 1711653199
transform 1 0 1116 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6212
timestamp 1711653199
transform 1 0 1092 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_6213
timestamp 1711653199
transform 1 0 1068 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6214
timestamp 1711653199
transform 1 0 1236 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6215
timestamp 1711653199
transform 1 0 1228 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6216
timestamp 1711653199
transform 1 0 1140 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6217
timestamp 1711653199
transform 1 0 1452 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6218
timestamp 1711653199
transform 1 0 1420 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6219
timestamp 1711653199
transform 1 0 1460 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6220
timestamp 1711653199
transform 1 0 1428 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6221
timestamp 1711653199
transform 1 0 1420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6222
timestamp 1711653199
transform 1 0 1060 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6223
timestamp 1711653199
transform 1 0 1692 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_6224
timestamp 1711653199
transform 1 0 1628 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_6225
timestamp 1711653199
transform 1 0 1628 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_6226
timestamp 1711653199
transform 1 0 1604 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_6227
timestamp 1711653199
transform 1 0 1468 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_6228
timestamp 1711653199
transform 1 0 1260 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6229
timestamp 1711653199
transform 1 0 1588 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6230
timestamp 1711653199
transform 1 0 1564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6231
timestamp 1711653199
transform 1 0 1596 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6232
timestamp 1711653199
transform 1 0 1532 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6233
timestamp 1711653199
transform 1 0 1516 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6234
timestamp 1711653199
transform 1 0 1108 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6235
timestamp 1711653199
transform 1 0 1772 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_6236
timestamp 1711653199
transform 1 0 1684 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6237
timestamp 1711653199
transform 1 0 1684 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6238
timestamp 1711653199
transform 1 0 1660 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6239
timestamp 1711653199
transform 1 0 1660 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6240
timestamp 1711653199
transform 1 0 1212 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6241
timestamp 1711653199
transform 1 0 1860 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6242
timestamp 1711653199
transform 1 0 1700 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6243
timestamp 1711653199
transform 1 0 1660 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6244
timestamp 1711653199
transform 1 0 1284 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6245
timestamp 1711653199
transform 1 0 1700 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_6246
timestamp 1711653199
transform 1 0 1292 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6247
timestamp 1711653199
transform 1 0 1236 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6248
timestamp 1711653199
transform 1 0 1164 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_6249
timestamp 1711653199
transform 1 0 1188 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_6250
timestamp 1711653199
transform 1 0 1172 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6251
timestamp 1711653199
transform 1 0 1284 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6252
timestamp 1711653199
transform 1 0 1260 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6253
timestamp 1711653199
transform 1 0 1228 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6254
timestamp 1711653199
transform 1 0 1164 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6255
timestamp 1711653199
transform 1 0 1316 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_6256
timestamp 1711653199
transform 1 0 1300 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6257
timestamp 1711653199
transform 1 0 1468 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_6258
timestamp 1711653199
transform 1 0 1284 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6259
timestamp 1711653199
transform 1 0 1180 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_6260
timestamp 1711653199
transform 1 0 1172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6261
timestamp 1711653199
transform 1 0 1724 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6262
timestamp 1711653199
transform 1 0 1692 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_6263
timestamp 1711653199
transform 1 0 1148 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6264
timestamp 1711653199
transform 1 0 1132 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6265
timestamp 1711653199
transform 1 0 732 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_6266
timestamp 1711653199
transform 1 0 724 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6267
timestamp 1711653199
transform 1 0 1948 0 1 2905
box -2 -2 2 2
use M2_M1  M2_M1_6268
timestamp 1711653199
transform 1 0 1932 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6269
timestamp 1711653199
transform 1 0 3212 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6270
timestamp 1711653199
transform 1 0 3180 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6271
timestamp 1711653199
transform 1 0 2740 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6272
timestamp 1711653199
transform 1 0 2652 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6273
timestamp 1711653199
transform 1 0 2060 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6274
timestamp 1711653199
transform 1 0 2044 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6275
timestamp 1711653199
transform 1 0 2404 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6276
timestamp 1711653199
transform 1 0 2388 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6277
timestamp 1711653199
transform 1 0 2516 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6278
timestamp 1711653199
transform 1 0 2508 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6279
timestamp 1711653199
transform 1 0 2188 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6280
timestamp 1711653199
transform 1 0 2140 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6281
timestamp 1711653199
transform 1 0 2244 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6282
timestamp 1711653199
transform 1 0 2228 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6283
timestamp 1711653199
transform 1 0 2548 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6284
timestamp 1711653199
transform 1 0 2460 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6285
timestamp 1711653199
transform 1 0 2468 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6286
timestamp 1711653199
transform 1 0 2412 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6287
timestamp 1711653199
transform 1 0 1972 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6288
timestamp 1711653199
transform 1 0 1940 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6289
timestamp 1711653199
transform 1 0 1844 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6290
timestamp 1711653199
transform 1 0 1812 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6291
timestamp 1711653199
transform 1 0 1612 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6292
timestamp 1711653199
transform 1 0 1580 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6293
timestamp 1711653199
transform 1 0 1724 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6294
timestamp 1711653199
transform 1 0 1708 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6295
timestamp 1711653199
transform 1 0 1492 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6296
timestamp 1711653199
transform 1 0 1444 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6297
timestamp 1711653199
transform 1 0 1332 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6298
timestamp 1711653199
transform 1 0 1332 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6299
timestamp 1711653199
transform 1 0 1068 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6300
timestamp 1711653199
transform 1 0 1068 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6301
timestamp 1711653199
transform 1 0 948 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6302
timestamp 1711653199
transform 1 0 924 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6303
timestamp 1711653199
transform 1 0 1188 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6304
timestamp 1711653199
transform 1 0 1188 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6305
timestamp 1711653199
transform 1 0 724 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6306
timestamp 1711653199
transform 1 0 628 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6307
timestamp 1711653199
transform 1 0 516 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6308
timestamp 1711653199
transform 1 0 516 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6309
timestamp 1711653199
transform 1 0 364 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6310
timestamp 1711653199
transform 1 0 364 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6311
timestamp 1711653199
transform 1 0 340 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6312
timestamp 1711653199
transform 1 0 300 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6313
timestamp 1711653199
transform 1 0 228 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6314
timestamp 1711653199
transform 1 0 220 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6315
timestamp 1711653199
transform 1 0 436 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6316
timestamp 1711653199
transform 1 0 356 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6317
timestamp 1711653199
transform 1 0 244 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6318
timestamp 1711653199
transform 1 0 140 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6319
timestamp 1711653199
transform 1 0 244 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6320
timestamp 1711653199
transform 1 0 132 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6321
timestamp 1711653199
transform 1 0 556 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6322
timestamp 1711653199
transform 1 0 468 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6323
timestamp 1711653199
transform 1 0 396 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6324
timestamp 1711653199
transform 1 0 324 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6325
timestamp 1711653199
transform 1 0 716 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6326
timestamp 1711653199
transform 1 0 604 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6327
timestamp 1711653199
transform 1 0 932 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6328
timestamp 1711653199
transform 1 0 836 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6329
timestamp 1711653199
transform 1 0 1412 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6330
timestamp 1711653199
transform 1 0 1316 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6331
timestamp 1711653199
transform 1 0 1588 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6332
timestamp 1711653199
transform 1 0 1548 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6333
timestamp 1711653199
transform 1 0 1772 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6334
timestamp 1711653199
transform 1 0 1764 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6335
timestamp 1711653199
transform 1 0 1908 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6336
timestamp 1711653199
transform 1 0 1868 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6337
timestamp 1711653199
transform 1 0 2988 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6338
timestamp 1711653199
transform 1 0 2852 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6339
timestamp 1711653199
transform 1 0 2852 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6340
timestamp 1711653199
transform 1 0 2948 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6341
timestamp 1711653199
transform 1 0 2948 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6342
timestamp 1711653199
transform 1 0 2940 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6343
timestamp 1711653199
transform 1 0 2940 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6344
timestamp 1711653199
transform 1 0 3004 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6345
timestamp 1711653199
transform 1 0 2956 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6346
timestamp 1711653199
transform 1 0 3036 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6347
timestamp 1711653199
transform 1 0 3004 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6348
timestamp 1711653199
transform 1 0 3340 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6349
timestamp 1711653199
transform 1 0 3300 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6350
timestamp 1711653199
transform 1 0 3028 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6351
timestamp 1711653199
transform 1 0 3020 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6352
timestamp 1711653199
transform 1 0 3356 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6353
timestamp 1711653199
transform 1 0 3252 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_6354
timestamp 1711653199
transform 1 0 3316 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6355
timestamp 1711653199
transform 1 0 3292 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6356
timestamp 1711653199
transform 1 0 3316 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6357
timestamp 1711653199
transform 1 0 3212 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6358
timestamp 1711653199
transform 1 0 3244 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6359
timestamp 1711653199
transform 1 0 3212 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6360
timestamp 1711653199
transform 1 0 3068 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6361
timestamp 1711653199
transform 1 0 3044 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6362
timestamp 1711653199
transform 1 0 3084 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6363
timestamp 1711653199
transform 1 0 3060 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6364
timestamp 1711653199
transform 1 0 3284 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6365
timestamp 1711653199
transform 1 0 3220 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6366
timestamp 1711653199
transform 1 0 3236 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6367
timestamp 1711653199
transform 1 0 3204 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6368
timestamp 1711653199
transform 1 0 3268 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6369
timestamp 1711653199
transform 1 0 3244 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6370
timestamp 1711653199
transform 1 0 3140 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6371
timestamp 1711653199
transform 1 0 3132 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6372
timestamp 1711653199
transform 1 0 3340 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6373
timestamp 1711653199
transform 1 0 3324 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6374
timestamp 1711653199
transform 1 0 3324 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_6375
timestamp 1711653199
transform 1 0 3140 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6376
timestamp 1711653199
transform 1 0 3092 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6377
timestamp 1711653199
transform 1 0 3084 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6378
timestamp 1711653199
transform 1 0 3068 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6379
timestamp 1711653199
transform 1 0 2988 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6380
timestamp 1711653199
transform 1 0 2980 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6381
timestamp 1711653199
transform 1 0 3220 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6382
timestamp 1711653199
transform 1 0 3116 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6383
timestamp 1711653199
transform 1 0 3100 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6384
timestamp 1711653199
transform 1 0 3132 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6385
timestamp 1711653199
transform 1 0 3116 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6386
timestamp 1711653199
transform 1 0 3196 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6387
timestamp 1711653199
transform 1 0 3004 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6388
timestamp 1711653199
transform 1 0 2988 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6389
timestamp 1711653199
transform 1 0 3028 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6390
timestamp 1711653199
transform 1 0 3004 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_6391
timestamp 1711653199
transform 1 0 3300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6392
timestamp 1711653199
transform 1 0 3228 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6393
timestamp 1711653199
transform 1 0 3100 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6394
timestamp 1711653199
transform 1 0 3036 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6395
timestamp 1711653199
transform 1 0 3028 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6396
timestamp 1711653199
transform 1 0 2852 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6397
timestamp 1711653199
transform 1 0 2828 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6398
timestamp 1711653199
transform 1 0 2796 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6399
timestamp 1711653199
transform 1 0 1620 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6400
timestamp 1711653199
transform 1 0 1596 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6401
timestamp 1711653199
transform 1 0 1380 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6402
timestamp 1711653199
transform 1 0 1348 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6403
timestamp 1711653199
transform 1 0 1340 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6404
timestamp 1711653199
transform 1 0 1092 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6405
timestamp 1711653199
transform 1 0 1060 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6406
timestamp 1711653199
transform 1 0 3060 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6407
timestamp 1711653199
transform 1 0 2676 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6408
timestamp 1711653199
transform 1 0 2572 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6409
timestamp 1711653199
transform 1 0 2388 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6410
timestamp 1711653199
transform 1 0 2340 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6411
timestamp 1711653199
transform 1 0 1924 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6412
timestamp 1711653199
transform 1 0 1908 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6413
timestamp 1711653199
transform 1 0 1884 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6414
timestamp 1711653199
transform 1 0 1604 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6415
timestamp 1711653199
transform 1 0 564 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6416
timestamp 1711653199
transform 1 0 492 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6417
timestamp 1711653199
transform 1 0 428 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6418
timestamp 1711653199
transform 1 0 188 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6419
timestamp 1711653199
transform 1 0 2268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6420
timestamp 1711653199
transform 1 0 2228 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6421
timestamp 1711653199
transform 1 0 1876 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6422
timestamp 1711653199
transform 1 0 1756 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6423
timestamp 1711653199
transform 1 0 1300 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6424
timestamp 1711653199
transform 1 0 1236 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6425
timestamp 1711653199
transform 1 0 2524 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6426
timestamp 1711653199
transform 1 0 2516 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_6427
timestamp 1711653199
transform 1 0 2516 0 1 1985
box -2 -2 2 2
use M2_M1  M2_M1_6428
timestamp 1711653199
transform 1 0 2284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6429
timestamp 1711653199
transform 1 0 1916 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6430
timestamp 1711653199
transform 1 0 1900 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6431
timestamp 1711653199
transform 1 0 1556 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6432
timestamp 1711653199
transform 1 0 1412 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6433
timestamp 1711653199
transform 1 0 2940 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6434
timestamp 1711653199
transform 1 0 2588 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6435
timestamp 1711653199
transform 1 0 2564 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6436
timestamp 1711653199
transform 1 0 2156 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6437
timestamp 1711653199
transform 1 0 1804 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6438
timestamp 1711653199
transform 1 0 1276 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6439
timestamp 1711653199
transform 1 0 2844 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6440
timestamp 1711653199
transform 1 0 2676 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6441
timestamp 1711653199
transform 1 0 2660 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6442
timestamp 1711653199
transform 1 0 2660 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6443
timestamp 1711653199
transform 1 0 1940 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6444
timestamp 1711653199
transform 1 0 1764 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6445
timestamp 1711653199
transform 1 0 1292 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6446
timestamp 1711653199
transform 1 0 2572 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6447
timestamp 1711653199
transform 1 0 2412 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6448
timestamp 1711653199
transform 1 0 2332 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6449
timestamp 1711653199
transform 1 0 2132 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6450
timestamp 1711653199
transform 1 0 1924 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6451
timestamp 1711653199
transform 1 0 1868 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6452
timestamp 1711653199
transform 1 0 1468 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6453
timestamp 1711653199
transform 1 0 2652 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6454
timestamp 1711653199
transform 1 0 2324 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6455
timestamp 1711653199
transform 1 0 2132 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6456
timestamp 1711653199
transform 1 0 2052 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6457
timestamp 1711653199
transform 1 0 1572 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6458
timestamp 1711653199
transform 1 0 2164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6459
timestamp 1711653199
transform 1 0 2132 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6460
timestamp 1711653199
transform 1 0 2124 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6461
timestamp 1711653199
transform 1 0 1652 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6462
timestamp 1711653199
transform 1 0 1644 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6463
timestamp 1711653199
transform 1 0 2092 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6464
timestamp 1711653199
transform 1 0 2060 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6465
timestamp 1711653199
transform 1 0 2028 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6466
timestamp 1711653199
transform 1 0 2020 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6467
timestamp 1711653199
transform 1 0 1748 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6468
timestamp 1711653199
transform 1 0 1708 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_6469
timestamp 1711653199
transform 1 0 2564 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6470
timestamp 1711653199
transform 1 0 2468 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6471
timestamp 1711653199
transform 1 0 2364 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6472
timestamp 1711653199
transform 1 0 2268 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6473
timestamp 1711653199
transform 1 0 2172 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6474
timestamp 1711653199
transform 1 0 2068 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6475
timestamp 1711653199
transform 1 0 1852 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6476
timestamp 1711653199
transform 1 0 2012 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6477
timestamp 1711653199
transform 1 0 1988 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6478
timestamp 1711653199
transform 1 0 1972 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6479
timestamp 1711653199
transform 1 0 1900 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6480
timestamp 1711653199
transform 1 0 1740 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6481
timestamp 1711653199
transform 1 0 1652 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6482
timestamp 1711653199
transform 1 0 1924 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6483
timestamp 1711653199
transform 1 0 1916 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6484
timestamp 1711653199
transform 1 0 1876 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6485
timestamp 1711653199
transform 1 0 1732 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_6486
timestamp 1711653199
transform 1 0 1724 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_6487
timestamp 1711653199
transform 1 0 1620 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6488
timestamp 1711653199
transform 1 0 1492 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6489
timestamp 1711653199
transform 1 0 1652 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6490
timestamp 1711653199
transform 1 0 1604 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6491
timestamp 1711653199
transform 1 0 1300 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6492
timestamp 1711653199
transform 1 0 1292 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6493
timestamp 1711653199
transform 1 0 1444 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6494
timestamp 1711653199
transform 1 0 1292 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6495
timestamp 1711653199
transform 1 0 1228 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6496
timestamp 1711653199
transform 1 0 1204 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6497
timestamp 1711653199
transform 1 0 1180 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6498
timestamp 1711653199
transform 1 0 1284 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6499
timestamp 1711653199
transform 1 0 1284 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6500
timestamp 1711653199
transform 1 0 1172 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6501
timestamp 1711653199
transform 1 0 1140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6502
timestamp 1711653199
transform 1 0 1140 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6503
timestamp 1711653199
transform 1 0 1124 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6504
timestamp 1711653199
transform 1 0 996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6505
timestamp 1711653199
transform 1 0 1140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6506
timestamp 1711653199
transform 1 0 1132 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_6507
timestamp 1711653199
transform 1 0 1124 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6508
timestamp 1711653199
transform 1 0 1108 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6509
timestamp 1711653199
transform 1 0 1100 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6510
timestamp 1711653199
transform 1 0 1076 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6511
timestamp 1711653199
transform 1 0 1012 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6512
timestamp 1711653199
transform 1 0 1268 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6513
timestamp 1711653199
transform 1 0 1132 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6514
timestamp 1711653199
transform 1 0 996 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6515
timestamp 1711653199
transform 1 0 876 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6516
timestamp 1711653199
transform 1 0 748 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6517
timestamp 1711653199
transform 1 0 348 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6518
timestamp 1711653199
transform 1 0 340 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6519
timestamp 1711653199
transform 1 0 1196 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6520
timestamp 1711653199
transform 1 0 1148 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6521
timestamp 1711653199
transform 1 0 732 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6522
timestamp 1711653199
transform 1 0 700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6523
timestamp 1711653199
transform 1 0 684 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6524
timestamp 1711653199
transform 1 0 516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_6525
timestamp 1711653199
transform 1 0 260 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6526
timestamp 1711653199
transform 1 0 236 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6527
timestamp 1711653199
transform 1 0 1084 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6528
timestamp 1711653199
transform 1 0 1076 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6529
timestamp 1711653199
transform 1 0 644 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6530
timestamp 1711653199
transform 1 0 636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6531
timestamp 1711653199
transform 1 0 268 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_6532
timestamp 1711653199
transform 1 0 220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6533
timestamp 1711653199
transform 1 0 212 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6534
timestamp 1711653199
transform 1 0 1044 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_6535
timestamp 1711653199
transform 1 0 1044 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_6536
timestamp 1711653199
transform 1 0 684 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6537
timestamp 1711653199
transform 1 0 676 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6538
timestamp 1711653199
transform 1 0 388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6539
timestamp 1711653199
transform 1 0 132 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6540
timestamp 1711653199
transform 1 0 100 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6541
timestamp 1711653199
transform 1 0 84 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_6542
timestamp 1711653199
transform 1 0 2676 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6543
timestamp 1711653199
transform 1 0 2676 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6544
timestamp 1711653199
transform 1 0 2452 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6545
timestamp 1711653199
transform 1 0 2388 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6546
timestamp 1711653199
transform 1 0 2380 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6547
timestamp 1711653199
transform 1 0 2140 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6548
timestamp 1711653199
transform 1 0 1788 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6549
timestamp 1711653199
transform 1 0 756 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6550
timestamp 1711653199
transform 1 0 604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_6551
timestamp 1711653199
transform 1 0 572 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6552
timestamp 1711653199
transform 1 0 532 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6553
timestamp 1711653199
transform 1 0 492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6554
timestamp 1711653199
transform 1 0 484 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6555
timestamp 1711653199
transform 1 0 700 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_6556
timestamp 1711653199
transform 1 0 604 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6557
timestamp 1711653199
transform 1 0 516 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6558
timestamp 1711653199
transform 1 0 516 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6559
timestamp 1711653199
transform 1 0 428 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6560
timestamp 1711653199
transform 1 0 420 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6561
timestamp 1711653199
transform 1 0 788 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6562
timestamp 1711653199
transform 1 0 756 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6563
timestamp 1711653199
transform 1 0 580 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6564
timestamp 1711653199
transform 1 0 556 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6565
timestamp 1711653199
transform 1 0 556 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6566
timestamp 1711653199
transform 1 0 540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6567
timestamp 1711653199
transform 1 0 540 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_6568
timestamp 1711653199
transform 1 0 988 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_6569
timestamp 1711653199
transform 1 0 972 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6570
timestamp 1711653199
transform 1 0 964 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6571
timestamp 1711653199
transform 1 0 876 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6572
timestamp 1711653199
transform 1 0 772 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_6573
timestamp 1711653199
transform 1 0 652 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6574
timestamp 1711653199
transform 1 0 644 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6575
timestamp 1711653199
transform 1 0 1220 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6576
timestamp 1711653199
transform 1 0 940 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6577
timestamp 1711653199
transform 1 0 924 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6578
timestamp 1711653199
transform 1 0 924 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6579
timestamp 1711653199
transform 1 0 764 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6580
timestamp 1711653199
transform 1 0 716 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6581
timestamp 1711653199
transform 1 0 988 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6582
timestamp 1711653199
transform 1 0 724 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6583
timestamp 1711653199
transform 1 0 660 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6584
timestamp 1711653199
transform 1 0 660 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6585
timestamp 1711653199
transform 1 0 636 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6586
timestamp 1711653199
transform 1 0 620 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6587
timestamp 1711653199
transform 1 0 1076 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6588
timestamp 1711653199
transform 1 0 812 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6589
timestamp 1711653199
transform 1 0 812 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6590
timestamp 1711653199
transform 1 0 724 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6591
timestamp 1711653199
transform 1 0 612 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6592
timestamp 1711653199
transform 1 0 604 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_6593
timestamp 1711653199
transform 1 0 572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6594
timestamp 1711653199
transform 1 0 1468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6595
timestamp 1711653199
transform 1 0 1428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6596
timestamp 1711653199
transform 1 0 1356 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6597
timestamp 1711653199
transform 1 0 1316 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6598
timestamp 1711653199
transform 1 0 876 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6599
timestamp 1711653199
transform 1 0 708 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_6600
timestamp 1711653199
transform 1 0 668 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6601
timestamp 1711653199
transform 1 0 1500 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6602
timestamp 1711653199
transform 1 0 1420 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6603
timestamp 1711653199
transform 1 0 1324 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6604
timestamp 1711653199
transform 1 0 1316 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_6605
timestamp 1711653199
transform 1 0 1308 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6606
timestamp 1711653199
transform 1 0 1308 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6607
timestamp 1711653199
transform 1 0 1164 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6608
timestamp 1711653199
transform 1 0 940 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6609
timestamp 1711653199
transform 1 0 1692 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6610
timestamp 1711653199
transform 1 0 1644 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6611
timestamp 1711653199
transform 1 0 1636 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6612
timestamp 1711653199
transform 1 0 1612 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_6613
timestamp 1711653199
transform 1 0 1428 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6614
timestamp 1711653199
transform 1 0 1148 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_6615
timestamp 1711653199
transform 1 0 956 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6616
timestamp 1711653199
transform 1 0 924 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6617
timestamp 1711653199
transform 1 0 2772 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_6618
timestamp 1711653199
transform 1 0 2420 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6619
timestamp 1711653199
transform 1 0 2084 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6620
timestamp 1711653199
transform 1 0 2068 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6621
timestamp 1711653199
transform 1 0 1980 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6622
timestamp 1711653199
transform 1 0 1892 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6623
timestamp 1711653199
transform 1 0 3212 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6624
timestamp 1711653199
transform 1 0 3156 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6625
timestamp 1711653199
transform 1 0 2884 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6626
timestamp 1711653199
transform 1 0 3124 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_6627
timestamp 1711653199
transform 1 0 1804 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_6628
timestamp 1711653199
transform 1 0 2100 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_6629
timestamp 1711653199
transform 1 0 2084 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6630
timestamp 1711653199
transform 1 0 2172 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6631
timestamp 1711653199
transform 1 0 2156 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6632
timestamp 1711653199
transform 1 0 2132 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6633
timestamp 1711653199
transform 1 0 2108 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6634
timestamp 1711653199
transform 1 0 2628 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6635
timestamp 1711653199
transform 1 0 2612 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6636
timestamp 1711653199
transform 1 0 2564 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6637
timestamp 1711653199
transform 1 0 2532 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6638
timestamp 1711653199
transform 1 0 2180 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6639
timestamp 1711653199
transform 1 0 2100 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6640
timestamp 1711653199
transform 1 0 2060 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6641
timestamp 1711653199
transform 1 0 2028 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6642
timestamp 1711653199
transform 1 0 2132 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6643
timestamp 1711653199
transform 1 0 2116 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6644
timestamp 1711653199
transform 1 0 2684 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6645
timestamp 1711653199
transform 1 0 2636 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6646
timestamp 1711653199
transform 1 0 2476 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6647
timestamp 1711653199
transform 1 0 2636 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6648
timestamp 1711653199
transform 1 0 2356 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6649
timestamp 1711653199
transform 1 0 2164 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6650
timestamp 1711653199
transform 1 0 1956 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6651
timestamp 1711653199
transform 1 0 2052 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_6652
timestamp 1711653199
transform 1 0 1956 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6653
timestamp 1711653199
transform 1 0 1924 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6654
timestamp 1711653199
transform 1 0 1236 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6655
timestamp 1711653199
transform 1 0 1124 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6656
timestamp 1711653199
transform 1 0 844 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6657
timestamp 1711653199
transform 1 0 1116 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_6658
timestamp 1711653199
transform 1 0 1092 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6659
timestamp 1711653199
transform 1 0 780 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6660
timestamp 1711653199
transform 1 0 900 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6661
timestamp 1711653199
transform 1 0 684 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6662
timestamp 1711653199
transform 1 0 948 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6663
timestamp 1711653199
transform 1 0 724 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6664
timestamp 1711653199
transform 1 0 740 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6665
timestamp 1711653199
transform 1 0 716 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6666
timestamp 1711653199
transform 1 0 700 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6667
timestamp 1711653199
transform 1 0 764 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_6668
timestamp 1711653199
transform 1 0 756 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_6669
timestamp 1711653199
transform 1 0 740 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_6670
timestamp 1711653199
transform 1 0 1036 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6671
timestamp 1711653199
transform 1 0 996 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6672
timestamp 1711653199
transform 1 0 820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6673
timestamp 1711653199
transform 1 0 780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6674
timestamp 1711653199
transform 1 0 860 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6675
timestamp 1711653199
transform 1 0 820 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6676
timestamp 1711653199
transform 1 0 756 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6677
timestamp 1711653199
transform 1 0 956 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6678
timestamp 1711653199
transform 1 0 804 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_6679
timestamp 1711653199
transform 1 0 764 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6680
timestamp 1711653199
transform 1 0 276 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_6681
timestamp 1711653199
transform 1 0 220 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_6682
timestamp 1711653199
transform 1 0 1148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6683
timestamp 1711653199
transform 1 0 1108 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6684
timestamp 1711653199
transform 1 0 1132 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6685
timestamp 1711653199
transform 1 0 1100 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6686
timestamp 1711653199
transform 1 0 1020 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6687
timestamp 1711653199
transform 1 0 1004 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6688
timestamp 1711653199
transform 1 0 972 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6689
timestamp 1711653199
transform 1 0 780 0 1 2595
box -2 -2 2 2
use M2_M1  M2_M1_6690
timestamp 1711653199
transform 1 0 1196 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6691
timestamp 1711653199
transform 1 0 1188 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_6692
timestamp 1711653199
transform 1 0 828 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6693
timestamp 1711653199
transform 1 0 1308 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6694
timestamp 1711653199
transform 1 0 1164 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_6695
timestamp 1711653199
transform 1 0 924 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_6696
timestamp 1711653199
transform 1 0 1708 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6697
timestamp 1711653199
transform 1 0 1684 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_6698
timestamp 1711653199
transform 1 0 3364 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_6699
timestamp 1711653199
transform 1 0 3348 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6700
timestamp 1711653199
transform 1 0 3292 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_6701
timestamp 1711653199
transform 1 0 3276 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_6702
timestamp 1711653199
transform 1 0 2468 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_6703
timestamp 1711653199
transform 1 0 2412 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6704
timestamp 1711653199
transform 1 0 2300 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6705
timestamp 1711653199
transform 1 0 2284 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6706
timestamp 1711653199
transform 1 0 2124 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6707
timestamp 1711653199
transform 1 0 1932 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6708
timestamp 1711653199
transform 1 0 1852 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6709
timestamp 1711653199
transform 1 0 1732 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6710
timestamp 1711653199
transform 1 0 1620 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6711
timestamp 1711653199
transform 1 0 1500 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6712
timestamp 1711653199
transform 1 0 1268 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6713
timestamp 1711653199
transform 1 0 1108 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6714
timestamp 1711653199
transform 1 0 956 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6715
timestamp 1711653199
transform 1 0 780 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_6716
timestamp 1711653199
transform 1 0 764 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_6717
timestamp 1711653199
transform 1 0 1788 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6718
timestamp 1711653199
transform 1 0 1764 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_6719
timestamp 1711653199
transform 1 0 2716 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6720
timestamp 1711653199
transform 1 0 2692 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6721
timestamp 1711653199
transform 1 0 2524 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_6722
timestamp 1711653199
transform 1 0 2492 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6723
timestamp 1711653199
transform 1 0 2340 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6724
timestamp 1711653199
transform 1 0 2220 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6725
timestamp 1711653199
transform 1 0 2092 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_6726
timestamp 1711653199
transform 1 0 1996 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1711653199
transform 1 0 2956 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1711653199
transform 1 0 2820 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1711653199
transform 1 0 2836 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1711653199
transform 1 0 2724 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1711653199
transform 1 0 2740 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1711653199
transform 1 0 2652 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1711653199
transform 1 0 2692 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1711653199
transform 1 0 2420 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1711653199
transform 1 0 2388 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1711653199
transform 1 0 2364 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1711653199
transform 1 0 2340 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1711653199
transform 1 0 2548 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1711653199
transform 1 0 2396 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1711653199
transform 1 0 2324 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_14
timestamp 1711653199
transform 1 0 2292 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1711653199
transform 1 0 2540 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1711653199
transform 1 0 2420 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1711653199
transform 1 0 2308 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1711653199
transform 1 0 2244 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1711653199
transform 1 0 2580 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1711653199
transform 1 0 2516 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1711653199
transform 1 0 2124 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1711653199
transform 1 0 2644 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1711653199
transform 1 0 2548 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1711653199
transform 1 0 2124 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1711653199
transform 1 0 2076 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1711653199
transform 1 0 3348 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1711653199
transform 1 0 3340 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1711653199
transform 1 0 3332 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1711653199
transform 1 0 3284 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1711653199
transform 1 0 2932 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1711653199
transform 1 0 2828 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1711653199
transform 1 0 2364 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1711653199
transform 1 0 2364 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1711653199
transform 1 0 2340 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1711653199
transform 1 0 2300 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1711653199
transform 1 0 1956 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1711653199
transform 1 0 1740 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1711653199
transform 1 0 1740 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1711653199
transform 1 0 948 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1711653199
transform 1 0 916 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1711653199
transform 1 0 900 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1711653199
transform 1 0 828 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1711653199
transform 1 0 828 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_44
timestamp 1711653199
transform 1 0 652 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1711653199
transform 1 0 604 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_46
timestamp 1711653199
transform 1 0 460 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1711653199
transform 1 0 460 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_48
timestamp 1711653199
transform 1 0 420 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_49
timestamp 1711653199
transform 1 0 420 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1711653199
transform 1 0 324 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_51
timestamp 1711653199
transform 1 0 268 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_52
timestamp 1711653199
transform 1 0 220 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1711653199
transform 1 0 84 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1711653199
transform 1 0 3060 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1711653199
transform 1 0 2916 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1711653199
transform 1 0 2884 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_57
timestamp 1711653199
transform 1 0 2828 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1711653199
transform 1 0 3404 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1711653199
transform 1 0 3404 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1711653199
transform 1 0 3116 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_61
timestamp 1711653199
transform 1 0 3004 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1711653199
transform 1 0 2980 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1711653199
transform 1 0 2924 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_64
timestamp 1711653199
transform 1 0 2828 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_65
timestamp 1711653199
transform 1 0 3020 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_66
timestamp 1711653199
transform 1 0 2980 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1711653199
transform 1 0 2980 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1711653199
transform 1 0 2964 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1711653199
transform 1 0 2956 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_70
timestamp 1711653199
transform 1 0 2948 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_71
timestamp 1711653199
transform 1 0 2892 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_72
timestamp 1711653199
transform 1 0 2892 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1711653199
transform 1 0 2836 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1711653199
transform 1 0 2788 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1711653199
transform 1 0 2772 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_76
timestamp 1711653199
transform 1 0 2740 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_77
timestamp 1711653199
transform 1 0 2724 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_78
timestamp 1711653199
transform 1 0 2884 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1711653199
transform 1 0 2860 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1711653199
transform 1 0 2836 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1711653199
transform 1 0 2836 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1711653199
transform 1 0 2804 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1711653199
transform 1 0 2804 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1711653199
transform 1 0 2796 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1711653199
transform 1 0 2788 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1711653199
transform 1 0 2756 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_87
timestamp 1711653199
transform 1 0 2716 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1711653199
transform 1 0 2692 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1711653199
transform 1 0 2660 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1711653199
transform 1 0 2636 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1711653199
transform 1 0 2724 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_92
timestamp 1711653199
transform 1 0 2692 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1711653199
transform 1 0 2684 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1711653199
transform 1 0 2684 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1711653199
transform 1 0 2652 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1711653199
transform 1 0 2620 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1711653199
transform 1 0 2620 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1711653199
transform 1 0 2596 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1711653199
transform 1 0 2596 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1711653199
transform 1 0 2588 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1711653199
transform 1 0 2572 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1711653199
transform 1 0 3372 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1711653199
transform 1 0 3204 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1711653199
transform 1 0 3124 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_105
timestamp 1711653199
transform 1 0 3116 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1711653199
transform 1 0 3100 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1711653199
transform 1 0 3092 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1711653199
transform 1 0 3068 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_109
timestamp 1711653199
transform 1 0 3068 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_110
timestamp 1711653199
transform 1 0 3300 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1711653199
transform 1 0 3300 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1711653199
transform 1 0 3196 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1711653199
transform 1 0 3108 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_114
timestamp 1711653199
transform 1 0 2076 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_115
timestamp 1711653199
transform 1 0 2020 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1711653199
transform 1 0 2572 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_117
timestamp 1711653199
transform 1 0 2468 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_118
timestamp 1711653199
transform 1 0 2604 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1711653199
transform 1 0 2508 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1711653199
transform 1 0 2476 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1711653199
transform 1 0 2380 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1711653199
transform 1 0 1980 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1711653199
transform 1 0 1916 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_124
timestamp 1711653199
transform 1 0 1740 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_125
timestamp 1711653199
transform 1 0 1684 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1711653199
transform 1 0 1372 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_127
timestamp 1711653199
transform 1 0 1276 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1711653199
transform 1 0 1100 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1711653199
transform 1 0 988 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1711653199
transform 1 0 956 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1711653199
transform 1 0 820 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1711653199
transform 1 0 1236 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1711653199
transform 1 0 1124 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1711653199
transform 1 0 548 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1711653199
transform 1 0 436 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1711653199
transform 1 0 396 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1711653199
transform 1 0 316 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1711653199
transform 1 0 396 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1711653199
transform 1 0 276 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1711653199
transform 1 0 252 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_141
timestamp 1711653199
transform 1 0 188 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1711653199
transform 1 0 396 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1711653199
transform 1 0 252 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1711653199
transform 1 0 3396 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1711653199
transform 1 0 3356 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1711653199
transform 1 0 3108 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1711653199
transform 1 0 2980 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1711653199
transform 1 0 2980 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1711653199
transform 1 0 2844 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1711653199
transform 1 0 2708 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1711653199
transform 1 0 2972 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1711653199
transform 1 0 2772 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1711653199
transform 1 0 2668 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1711653199
transform 1 0 2316 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1711653199
transform 1 0 1964 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1711653199
transform 1 0 2412 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1711653199
transform 1 0 2372 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1711653199
transform 1 0 2380 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1711653199
transform 1 0 2156 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1711653199
transform 1 0 2268 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1711653199
transform 1 0 2116 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1711653199
transform 1 0 2524 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1711653199
transform 1 0 2308 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1711653199
transform 1 0 2636 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1711653199
transform 1 0 2548 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1711653199
transform 1 0 2116 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1711653199
transform 1 0 1900 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1711653199
transform 1 0 2276 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1711653199
transform 1 0 1868 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1711653199
transform 1 0 1708 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1711653199
transform 1 0 1628 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1711653199
transform 1 0 1484 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1711653199
transform 1 0 1348 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1711653199
transform 1 0 660 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1711653199
transform 1 0 596 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1711653199
transform 1 0 508 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1711653199
transform 1 0 388 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1711653199
transform 1 0 524 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1711653199
transform 1 0 460 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1711653199
transform 1 0 380 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_181
timestamp 1711653199
transform 1 0 332 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1711653199
transform 1 0 1124 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1711653199
transform 1 0 1092 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1711653199
transform 1 0 1236 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1711653199
transform 1 0 1124 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_186
timestamp 1711653199
transform 1 0 1436 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1711653199
transform 1 0 1188 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1711653199
transform 1 0 1596 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1711653199
transform 1 0 1276 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1711653199
transform 1 0 1868 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1711653199
transform 1 0 1604 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1711653199
transform 1 0 2012 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1711653199
transform 1 0 1884 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1711653199
transform 1 0 2116 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1711653199
transform 1 0 2076 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1711653199
transform 1 0 2220 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1711653199
transform 1 0 2124 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1711653199
transform 1 0 2796 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1711653199
transform 1 0 2700 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1711653199
transform 1 0 1788 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1711653199
transform 1 0 1660 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1711653199
transform 1 0 1548 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1711653199
transform 1 0 1452 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1711653199
transform 1 0 1084 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1711653199
transform 1 0 988 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1711653199
transform 1 0 908 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1711653199
transform 1 0 780 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1711653199
transform 1 0 572 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1711653199
transform 1 0 508 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1711653199
transform 1 0 500 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_211
timestamp 1711653199
transform 1 0 364 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1711653199
transform 1 0 284 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1711653199
transform 1 0 196 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1711653199
transform 1 0 1116 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1711653199
transform 1 0 508 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1711653199
transform 1 0 1164 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1711653199
transform 1 0 436 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1711653199
transform 1 0 1220 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1711653199
transform 1 0 828 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1711653199
transform 1 0 1316 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1711653199
transform 1 0 1076 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1711653199
transform 1 0 2100 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1711653199
transform 1 0 1932 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1711653199
transform 1 0 2148 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1711653199
transform 1 0 2068 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1711653199
transform 1 0 3212 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1711653199
transform 1 0 3212 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_228
timestamp 1711653199
transform 1 0 3180 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1711653199
transform 1 0 3052 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1711653199
transform 1 0 3020 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1711653199
transform 1 0 2924 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1711653199
transform 1 0 2660 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1711653199
transform 1 0 3276 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1711653199
transform 1 0 3252 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1711653199
transform 1 0 3220 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_236
timestamp 1711653199
transform 1 0 3220 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1711653199
transform 1 0 3044 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1711653199
transform 1 0 3044 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1711653199
transform 1 0 2996 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1711653199
transform 1 0 2940 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_241
timestamp 1711653199
transform 1 0 2516 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1711653199
transform 1 0 2844 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_243
timestamp 1711653199
transform 1 0 2500 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_244
timestamp 1711653199
transform 1 0 2812 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_245
timestamp 1711653199
transform 1 0 2788 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_246
timestamp 1711653199
transform 1 0 2772 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1711653199
transform 1 0 2716 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_248
timestamp 1711653199
transform 1 0 2548 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1711653199
transform 1 0 2868 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1711653199
transform 1 0 2740 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_251
timestamp 1711653199
transform 1 0 2684 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1711653199
transform 1 0 2684 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_253
timestamp 1711653199
transform 1 0 2612 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1711653199
transform 1 0 3380 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1711653199
transform 1 0 3356 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1711653199
transform 1 0 3316 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1711653199
transform 1 0 3164 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_258
timestamp 1711653199
transform 1 0 3124 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_259
timestamp 1711653199
transform 1 0 3028 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1711653199
transform 1 0 3324 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1711653199
transform 1 0 3292 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1711653199
transform 1 0 3252 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1711653199
transform 1 0 3212 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_264
timestamp 1711653199
transform 1 0 3348 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_265
timestamp 1711653199
transform 1 0 3260 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_266
timestamp 1711653199
transform 1 0 3260 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1711653199
transform 1 0 3204 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_268
timestamp 1711653199
transform 1 0 3196 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_269
timestamp 1711653199
transform 1 0 3188 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1711653199
transform 1 0 3164 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_271
timestamp 1711653199
transform 1 0 3156 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_272
timestamp 1711653199
transform 1 0 3148 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1711653199
transform 1 0 3020 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_274
timestamp 1711653199
transform 1 0 2948 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1711653199
transform 1 0 2820 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1711653199
transform 1 0 2924 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_277
timestamp 1711653199
transform 1 0 2788 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_278
timestamp 1711653199
transform 1 0 2956 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1711653199
transform 1 0 2844 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_280
timestamp 1711653199
transform 1 0 3396 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_281
timestamp 1711653199
transform 1 0 3300 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1711653199
transform 1 0 3260 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1711653199
transform 1 0 3260 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1711653199
transform 1 0 3228 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1711653199
transform 1 0 3156 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_286
timestamp 1711653199
transform 1 0 3140 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_287
timestamp 1711653199
transform 1 0 3084 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1711653199
transform 1 0 3028 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1711653199
transform 1 0 3220 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_290
timestamp 1711653199
transform 1 0 3132 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1711653199
transform 1 0 3100 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1711653199
transform 1 0 3388 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1711653199
transform 1 0 3244 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1711653199
transform 1 0 3172 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1711653199
transform 1 0 3172 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1711653199
transform 1 0 3084 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1711653199
transform 1 0 3076 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1711653199
transform 1 0 3060 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1711653199
transform 1 0 3052 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1711653199
transform 1 0 2964 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1711653199
transform 1 0 2836 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1711653199
transform 1 0 2740 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1711653199
transform 1 0 3044 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1711653199
transform 1 0 2980 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1711653199
transform 1 0 3236 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1711653199
transform 1 0 3236 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1711653199
transform 1 0 3220 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1711653199
transform 1 0 3212 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1711653199
transform 1 0 3212 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_310
timestamp 1711653199
transform 1 0 3204 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1711653199
transform 1 0 3164 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1711653199
transform 1 0 3124 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1711653199
transform 1 0 2916 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1711653199
transform 1 0 2772 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1711653199
transform 1 0 2756 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1711653199
transform 1 0 3260 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1711653199
transform 1 0 3260 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1711653199
transform 1 0 3236 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1711653199
transform 1 0 3180 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1711653199
transform 1 0 3132 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1711653199
transform 1 0 3252 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1711653199
transform 1 0 3044 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_323
timestamp 1711653199
transform 1 0 2212 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1711653199
transform 1 0 2124 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1711653199
transform 1 0 2124 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1711653199
transform 1 0 2028 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1711653199
transform 1 0 1892 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_328
timestamp 1711653199
transform 1 0 1876 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1711653199
transform 1 0 1660 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1711653199
transform 1 0 1628 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1711653199
transform 1 0 1564 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1711653199
transform 1 0 1500 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1711653199
transform 1 0 1492 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1711653199
transform 1 0 844 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1711653199
transform 1 0 844 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1711653199
transform 1 0 772 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1711653199
transform 1 0 540 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1711653199
transform 1 0 468 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_339
timestamp 1711653199
transform 1 0 468 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_340
timestamp 1711653199
transform 1 0 380 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1711653199
transform 1 0 372 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1711653199
transform 1 0 292 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1711653199
transform 1 0 292 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1711653199
transform 1 0 268 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1711653199
transform 1 0 268 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1711653199
transform 1 0 244 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1711653199
transform 1 0 244 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1711653199
transform 1 0 3044 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_349
timestamp 1711653199
transform 1 0 3036 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1711653199
transform 1 0 2836 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1711653199
transform 1 0 2660 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_352
timestamp 1711653199
transform 1 0 2652 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_353
timestamp 1711653199
transform 1 0 2612 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1711653199
transform 1 0 2580 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_355
timestamp 1711653199
transform 1 0 2476 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1711653199
transform 1 0 2476 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1711653199
transform 1 0 2452 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1711653199
transform 1 0 2380 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1711653199
transform 1 0 2364 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_360
timestamp 1711653199
transform 1 0 2348 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1711653199
transform 1 0 2180 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1711653199
transform 1 0 2180 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1711653199
transform 1 0 2164 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1711653199
transform 1 0 1876 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_365
timestamp 1711653199
transform 1 0 1876 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_366
timestamp 1711653199
transform 1 0 1828 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1711653199
transform 1 0 1788 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1711653199
transform 1 0 1780 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1711653199
transform 1 0 1172 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1711653199
transform 1 0 1172 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1711653199
transform 1 0 956 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1711653199
transform 1 0 948 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1711653199
transform 1 0 908 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1711653199
transform 1 0 908 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1711653199
transform 1 0 716 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1711653199
transform 1 0 716 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1711653199
transform 1 0 668 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1711653199
transform 1 0 1532 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1711653199
transform 1 0 1260 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1711653199
transform 1 0 1084 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_381
timestamp 1711653199
transform 1 0 2892 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1711653199
transform 1 0 2892 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1711653199
transform 1 0 2828 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1711653199
transform 1 0 2812 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1711653199
transform 1 0 2796 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1711653199
transform 1 0 2788 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1711653199
transform 1 0 2788 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1711653199
transform 1 0 2756 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1711653199
transform 1 0 2748 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_390
timestamp 1711653199
transform 1 0 2748 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1711653199
transform 1 0 2676 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1711653199
transform 1 0 2676 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1711653199
transform 1 0 1716 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_394
timestamp 1711653199
transform 1 0 1692 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1711653199
transform 1 0 1652 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1711653199
transform 1 0 2852 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1711653199
transform 1 0 2772 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1711653199
transform 1 0 2684 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1711653199
transform 1 0 2988 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1711653199
transform 1 0 2940 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1711653199
transform 1 0 2892 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1711653199
transform 1 0 2892 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1711653199
transform 1 0 2836 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1711653199
transform 1 0 2836 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1711653199
transform 1 0 2812 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1711653199
transform 1 0 2804 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1711653199
transform 1 0 2804 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1711653199
transform 1 0 2772 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1711653199
transform 1 0 2740 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1711653199
transform 1 0 2740 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1711653199
transform 1 0 2716 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_412
timestamp 1711653199
transform 1 0 2652 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1711653199
transform 1 0 2308 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1711653199
transform 1 0 2308 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_415
timestamp 1711653199
transform 1 0 1324 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1711653199
transform 1 0 2612 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1711653199
transform 1 0 2548 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1711653199
transform 1 0 2492 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1711653199
transform 1 0 2436 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1711653199
transform 1 0 2420 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_421
timestamp 1711653199
transform 1 0 2340 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1711653199
transform 1 0 2300 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1711653199
transform 1 0 2220 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1711653199
transform 1 0 2212 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1711653199
transform 1 0 2204 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1711653199
transform 1 0 2028 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1711653199
transform 1 0 972 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1711653199
transform 1 0 972 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1711653199
transform 1 0 884 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1711653199
transform 1 0 884 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1711653199
transform 1 0 516 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1711653199
transform 1 0 516 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1711653199
transform 1 0 356 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1711653199
transform 1 0 332 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1711653199
transform 1 0 212 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1711653199
transform 1 0 196 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1711653199
transform 1 0 1788 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1711653199
transform 1 0 1724 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1711653199
transform 1 0 1724 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1711653199
transform 1 0 1548 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1711653199
transform 1 0 1524 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1711653199
transform 1 0 1476 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1711653199
transform 1 0 1380 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1711653199
transform 1 0 1380 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1711653199
transform 1 0 1316 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1711653199
transform 1 0 2964 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1711653199
transform 1 0 2964 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1711653199
transform 1 0 2956 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1711653199
transform 1 0 2932 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1711653199
transform 1 0 2924 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1711653199
transform 1 0 2876 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1711653199
transform 1 0 2868 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1711653199
transform 1 0 2812 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1711653199
transform 1 0 2284 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1711653199
transform 1 0 2252 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1711653199
transform 1 0 2948 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1711653199
transform 1 0 2892 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1711653199
transform 1 0 2884 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1711653199
transform 1 0 2852 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1711653199
transform 1 0 740 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1711653199
transform 1 0 732 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1711653199
transform 1 0 708 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1711653199
transform 1 0 708 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1711653199
transform 1 0 700 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1711653199
transform 1 0 700 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1711653199
transform 1 0 700 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1711653199
transform 1 0 676 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1711653199
transform 1 0 668 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1711653199
transform 1 0 668 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1711653199
transform 1 0 516 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1711653199
transform 1 0 508 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1711653199
transform 1 0 508 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1711653199
transform 1 0 428 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1711653199
transform 1 0 3404 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_475
timestamp 1711653199
transform 1 0 3340 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1711653199
transform 1 0 3044 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1711653199
transform 1 0 1468 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_478
timestamp 1711653199
transform 1 0 1172 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1711653199
transform 1 0 1052 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1711653199
transform 1 0 1052 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1711653199
transform 1 0 636 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1711653199
transform 1 0 636 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1711653199
transform 1 0 636 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1711653199
transform 1 0 612 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1711653199
transform 1 0 612 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1711653199
transform 1 0 596 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1711653199
transform 1 0 572 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1711653199
transform 1 0 548 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_489
timestamp 1711653199
transform 1 0 484 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1711653199
transform 1 0 484 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1711653199
transform 1 0 484 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1711653199
transform 1 0 92 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1711653199
transform 1 0 3236 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1711653199
transform 1 0 3228 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1711653199
transform 1 0 3180 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1711653199
transform 1 0 3132 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1711653199
transform 1 0 3044 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1711653199
transform 1 0 3044 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1711653199
transform 1 0 2588 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_500
timestamp 1711653199
transform 1 0 2588 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1711653199
transform 1 0 2516 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1711653199
transform 1 0 2468 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_503
timestamp 1711653199
transform 1 0 2452 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_504
timestamp 1711653199
transform 1 0 2364 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_505
timestamp 1711653199
transform 1 0 2356 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_506
timestamp 1711653199
transform 1 0 2044 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_507
timestamp 1711653199
transform 1 0 2036 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1711653199
transform 1 0 1996 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1711653199
transform 1 0 1988 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1711653199
transform 1 0 1988 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1711653199
transform 1 0 1908 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1711653199
transform 1 0 1348 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_513
timestamp 1711653199
transform 1 0 1324 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1711653199
transform 1 0 1324 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1711653199
transform 1 0 716 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_516
timestamp 1711653199
transform 1 0 700 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_517
timestamp 1711653199
transform 1 0 700 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1711653199
transform 1 0 700 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1711653199
transform 1 0 700 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1711653199
transform 1 0 604 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1711653199
transform 1 0 604 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1711653199
transform 1 0 572 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1711653199
transform 1 0 572 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1711653199
transform 1 0 564 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_525
timestamp 1711653199
transform 1 0 556 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1711653199
transform 1 0 500 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_527
timestamp 1711653199
transform 1 0 492 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1711653199
transform 1 0 1228 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1711653199
transform 1 0 1164 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1711653199
transform 1 0 876 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1711653199
transform 1 0 876 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_532
timestamp 1711653199
transform 1 0 844 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_533
timestamp 1711653199
transform 1 0 804 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1711653199
transform 1 0 804 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1711653199
transform 1 0 748 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_536
timestamp 1711653199
transform 1 0 740 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_537
timestamp 1711653199
transform 1 0 724 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1711653199
transform 1 0 3052 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_539
timestamp 1711653199
transform 1 0 2964 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_540
timestamp 1711653199
transform 1 0 2956 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_541
timestamp 1711653199
transform 1 0 2940 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_542
timestamp 1711653199
transform 1 0 2924 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_543
timestamp 1711653199
transform 1 0 2908 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1711653199
transform 1 0 2908 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_545
timestamp 1711653199
transform 1 0 2908 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_546
timestamp 1711653199
transform 1 0 1396 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1711653199
transform 1 0 2204 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1711653199
transform 1 0 2180 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_549
timestamp 1711653199
transform 1 0 2092 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1711653199
transform 1 0 1940 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1711653199
transform 1 0 1836 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1711653199
transform 1 0 2172 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_553
timestamp 1711653199
transform 1 0 2156 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1711653199
transform 1 0 2148 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1711653199
transform 1 0 2116 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_556
timestamp 1711653199
transform 1 0 2116 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_557
timestamp 1711653199
transform 1 0 1980 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_558
timestamp 1711653199
transform 1 0 1956 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1711653199
transform 1 0 652 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_560
timestamp 1711653199
transform 1 0 620 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_561
timestamp 1711653199
transform 1 0 620 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_562
timestamp 1711653199
transform 1 0 420 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1711653199
transform 1 0 228 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1711653199
transform 1 0 228 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1711653199
transform 1 0 180 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1711653199
transform 1 0 180 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_567
timestamp 1711653199
transform 1 0 156 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1711653199
transform 1 0 156 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_569
timestamp 1711653199
transform 1 0 156 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1711653199
transform 1 0 132 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_571
timestamp 1711653199
transform 1 0 108 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1711653199
transform 1 0 108 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_573
timestamp 1711653199
transform 1 0 2236 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1711653199
transform 1 0 2132 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1711653199
transform 1 0 2132 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1711653199
transform 1 0 2044 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1711653199
transform 1 0 2044 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1711653199
transform 1 0 1852 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1711653199
transform 1 0 1820 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1711653199
transform 1 0 1812 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1711653199
transform 1 0 1804 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1711653199
transform 1 0 1524 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1711653199
transform 1 0 1364 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1711653199
transform 1 0 1364 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1711653199
transform 1 0 956 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1711653199
transform 1 0 276 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_587
timestamp 1711653199
transform 1 0 260 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1711653199
transform 1 0 196 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1711653199
transform 1 0 3356 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1711653199
transform 1 0 3332 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1711653199
transform 1 0 3108 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1711653199
transform 1 0 2996 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1711653199
transform 1 0 2996 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1711653199
transform 1 0 2940 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1711653199
transform 1 0 2940 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_596
timestamp 1711653199
transform 1 0 2588 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1711653199
transform 1 0 2532 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1711653199
transform 1 0 2532 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1711653199
transform 1 0 2452 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1711653199
transform 1 0 2452 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1711653199
transform 1 0 1908 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1711653199
transform 1 0 3116 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1711653199
transform 1 0 2804 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1711653199
transform 1 0 2684 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1711653199
transform 1 0 2316 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_606
timestamp 1711653199
transform 1 0 1580 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1711653199
transform 1 0 1580 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1711653199
transform 1 0 1084 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1711653199
transform 1 0 1044 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1711653199
transform 1 0 1028 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1711653199
transform 1 0 1028 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1711653199
transform 1 0 1028 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1711653199
transform 1 0 2940 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1711653199
transform 1 0 2932 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1711653199
transform 1 0 2884 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1711653199
transform 1 0 2876 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_617
timestamp 1711653199
transform 1 0 2836 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1711653199
transform 1 0 2828 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1711653199
transform 1 0 2812 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1711653199
transform 1 0 2796 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1711653199
transform 1 0 2780 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1711653199
transform 1 0 2764 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1711653199
transform 1 0 2580 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1711653199
transform 1 0 2580 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1711653199
transform 1 0 2524 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1711653199
transform 1 0 2524 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1711653199
transform 1 0 2236 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1711653199
transform 1 0 2236 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1711653199
transform 1 0 2020 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1711653199
transform 1 0 2620 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1711653199
transform 1 0 2596 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1711653199
transform 1 0 2588 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1711653199
transform 1 0 2588 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1711653199
transform 1 0 2556 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1711653199
transform 1 0 2540 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1711653199
transform 1 0 2260 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1711653199
transform 1 0 316 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1711653199
transform 1 0 2140 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1711653199
transform 1 0 2140 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1711653199
transform 1 0 2140 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1711653199
transform 1 0 2108 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1711653199
transform 1 0 2100 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_643
timestamp 1711653199
transform 1 0 2084 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1711653199
transform 1 0 2100 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1711653199
transform 1 0 2076 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1711653199
transform 1 0 1900 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1711653199
transform 1 0 1596 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1711653199
transform 1 0 1596 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1711653199
transform 1 0 1204 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1711653199
transform 1 0 1204 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1711653199
transform 1 0 1076 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1711653199
transform 1 0 756 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_653
timestamp 1711653199
transform 1 0 756 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_654
timestamp 1711653199
transform 1 0 500 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1711653199
transform 1 0 436 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1711653199
transform 1 0 2756 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1711653199
transform 1 0 2724 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1711653199
transform 1 0 2724 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1711653199
transform 1 0 2676 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1711653199
transform 1 0 2604 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1711653199
transform 1 0 2532 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1711653199
transform 1 0 2252 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1711653199
transform 1 0 2236 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1711653199
transform 1 0 2212 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1711653199
transform 1 0 1548 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1711653199
transform 1 0 2612 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1711653199
transform 1 0 2556 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1711653199
transform 1 0 1012 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1711653199
transform 1 0 1004 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1711653199
transform 1 0 940 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1711653199
transform 1 0 932 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1711653199
transform 1 0 860 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1711653199
transform 1 0 2668 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1711653199
transform 1 0 2660 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1711653199
transform 1 0 2308 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_676
timestamp 1711653199
transform 1 0 2308 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_677
timestamp 1711653199
transform 1 0 2292 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1711653199
transform 1 0 2076 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1711653199
transform 1 0 2076 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1711653199
transform 1 0 2044 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1711653199
transform 1 0 2020 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1711653199
transform 1 0 1380 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1711653199
transform 1 0 1380 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1711653199
transform 1 0 1372 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1711653199
transform 1 0 1212 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1711653199
transform 1 0 1204 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1711653199
transform 1 0 1148 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1711653199
transform 1 0 1140 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1711653199
transform 1 0 836 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1711653199
transform 1 0 836 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1711653199
transform 1 0 452 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1711653199
transform 1 0 444 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_693
timestamp 1711653199
transform 1 0 388 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1711653199
transform 1 0 380 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1711653199
transform 1 0 340 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1711653199
transform 1 0 340 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1711653199
transform 1 0 588 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1711653199
transform 1 0 588 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1711653199
transform 1 0 588 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1711653199
transform 1 0 588 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1711653199
transform 1 0 564 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1711653199
transform 1 0 556 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1711653199
transform 1 0 556 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1711653199
transform 1 0 532 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1711653199
transform 1 0 532 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_706
timestamp 1711653199
transform 1 0 516 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_707
timestamp 1711653199
transform 1 0 484 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1711653199
transform 1 0 476 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1711653199
transform 1 0 468 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1711653199
transform 1 0 468 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1711653199
transform 1 0 444 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1711653199
transform 1 0 436 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1711653199
transform 1 0 348 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1711653199
transform 1 0 348 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1711653199
transform 1 0 252 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1711653199
transform 1 0 228 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_717
timestamp 1711653199
transform 1 0 156 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1711653199
transform 1 0 148 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_719
timestamp 1711653199
transform 1 0 108 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1711653199
transform 1 0 3372 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1711653199
transform 1 0 3372 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1711653199
transform 1 0 3356 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1711653199
transform 1 0 3356 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1711653199
transform 1 0 3332 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1711653199
transform 1 0 3316 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1711653199
transform 1 0 1396 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_727
timestamp 1711653199
transform 1 0 1396 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1711653199
transform 1 0 1364 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1711653199
transform 1 0 1364 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1711653199
transform 1 0 1364 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1711653199
transform 1 0 1364 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1711653199
transform 1 0 1316 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1711653199
transform 1 0 1316 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1711653199
transform 1 0 1300 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1711653199
transform 1 0 1276 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1711653199
transform 1 0 1244 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1711653199
transform 1 0 1204 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1711653199
transform 1 0 1140 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1711653199
transform 1 0 1140 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1711653199
transform 1 0 3196 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1711653199
transform 1 0 3196 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1711653199
transform 1 0 3116 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1711653199
transform 1 0 3108 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1711653199
transform 1 0 3092 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1711653199
transform 1 0 3092 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1711653199
transform 1 0 3052 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1711653199
transform 1 0 2612 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1711653199
transform 1 0 2612 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1711653199
transform 1 0 2556 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1711653199
transform 1 0 2556 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1711653199
transform 1 0 2524 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1711653199
transform 1 0 2300 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1711653199
transform 1 0 2284 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1711653199
transform 1 0 3324 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1711653199
transform 1 0 3316 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1711653199
transform 1 0 3308 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1711653199
transform 1 0 3308 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1711653199
transform 1 0 3292 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1711653199
transform 1 0 3284 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1711653199
transform 1 0 3268 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1711653199
transform 1 0 2412 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1711653199
transform 1 0 2372 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1711653199
transform 1 0 2372 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1711653199
transform 1 0 2212 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1711653199
transform 1 0 364 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1711653199
transform 1 0 364 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_767
timestamp 1711653199
transform 1 0 356 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1711653199
transform 1 0 356 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1711653199
transform 1 0 332 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1711653199
transform 1 0 316 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1711653199
transform 1 0 316 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1711653199
transform 1 0 308 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1711653199
transform 1 0 308 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1711653199
transform 1 0 308 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1711653199
transform 1 0 300 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1711653199
transform 1 0 284 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1711653199
transform 1 0 276 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1711653199
transform 1 0 268 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1711653199
transform 1 0 268 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1711653199
transform 1 0 220 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1711653199
transform 1 0 212 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1711653199
transform 1 0 212 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1711653199
transform 1 0 180 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1711653199
transform 1 0 180 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1711653199
transform 1 0 3364 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1711653199
transform 1 0 3364 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1711653199
transform 1 0 3340 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_788
timestamp 1711653199
transform 1 0 3340 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1711653199
transform 1 0 3300 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1711653199
transform 1 0 3292 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1711653199
transform 1 0 3180 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_792
timestamp 1711653199
transform 1 0 3140 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1711653199
transform 1 0 3140 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1711653199
transform 1 0 2604 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1711653199
transform 1 0 2604 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1711653199
transform 1 0 2348 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_797
timestamp 1711653199
transform 1 0 2348 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1711653199
transform 1 0 2148 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1711653199
transform 1 0 356 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1711653199
transform 1 0 340 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1711653199
transform 1 0 340 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1711653199
transform 1 0 324 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_803
timestamp 1711653199
transform 1 0 324 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1711653199
transform 1 0 316 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_805
timestamp 1711653199
transform 1 0 316 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1711653199
transform 1 0 308 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1711653199
transform 1 0 308 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_808
timestamp 1711653199
transform 1 0 308 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1711653199
transform 1 0 300 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1711653199
transform 1 0 300 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1711653199
transform 1 0 292 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1711653199
transform 1 0 292 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1711653199
transform 1 0 276 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1711653199
transform 1 0 276 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1711653199
transform 1 0 260 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_816
timestamp 1711653199
transform 1 0 236 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1711653199
transform 1 0 236 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1711653199
transform 1 0 196 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1711653199
transform 1 0 188 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1711653199
transform 1 0 188 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1711653199
transform 1 0 116 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_822
timestamp 1711653199
transform 1 0 108 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1711653199
transform 1 0 2180 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1711653199
transform 1 0 2156 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1711653199
transform 1 0 2156 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1711653199
transform 1 0 2044 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1711653199
transform 1 0 1852 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1711653199
transform 1 0 1412 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1711653199
transform 1 0 1372 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1711653199
transform 1 0 1324 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1711653199
transform 1 0 628 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1711653199
transform 1 0 620 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1711653199
transform 1 0 572 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1711653199
transform 1 0 572 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_835
timestamp 1711653199
transform 1 0 428 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1711653199
transform 1 0 428 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1711653199
transform 1 0 308 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1711653199
transform 1 0 268 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1711653199
transform 1 0 268 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_840
timestamp 1711653199
transform 1 0 236 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1711653199
transform 1 0 196 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_842
timestamp 1711653199
transform 1 0 196 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1711653199
transform 1 0 1164 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1711653199
transform 1 0 1084 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_845
timestamp 1711653199
transform 1 0 1020 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1711653199
transform 1 0 1020 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_847
timestamp 1711653199
transform 1 0 820 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1711653199
transform 1 0 620 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1711653199
transform 1 0 476 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1711653199
transform 1 0 476 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1711653199
transform 1 0 452 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1711653199
transform 1 0 436 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1711653199
transform 1 0 388 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1711653199
transform 1 0 3356 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1711653199
transform 1 0 3252 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1711653199
transform 1 0 2908 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_857
timestamp 1711653199
transform 1 0 2900 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1711653199
transform 1 0 2876 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1711653199
transform 1 0 2860 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_860
timestamp 1711653199
transform 1 0 2860 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1711653199
transform 1 0 2772 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1711653199
transform 1 0 2772 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1711653199
transform 1 0 2540 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1711653199
transform 1 0 2540 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1711653199
transform 1 0 1348 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_866
timestamp 1711653199
transform 1 0 2612 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1711653199
transform 1 0 2612 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1711653199
transform 1 0 2580 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1711653199
transform 1 0 2580 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1711653199
transform 1 0 2244 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1711653199
transform 1 0 2172 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_872
timestamp 1711653199
transform 1 0 2172 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1711653199
transform 1 0 2108 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_874
timestamp 1711653199
transform 1 0 2100 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1711653199
transform 1 0 2092 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1711653199
transform 1 0 2092 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1711653199
transform 1 0 2028 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1711653199
transform 1 0 1700 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1711653199
transform 1 0 1252 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1711653199
transform 1 0 1220 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1711653199
transform 1 0 1220 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1711653199
transform 1 0 1156 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1711653199
transform 1 0 588 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1711653199
transform 1 0 588 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1711653199
transform 1 0 532 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1711653199
transform 1 0 532 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1711653199
transform 1 0 532 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1711653199
transform 1 0 484 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1711653199
transform 1 0 420 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1711653199
transform 1 0 420 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1711653199
transform 1 0 388 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1711653199
transform 1 0 388 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1711653199
transform 1 0 252 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1711653199
transform 1 0 252 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1711653199
transform 1 0 2204 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1711653199
transform 1 0 2204 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1711653199
transform 1 0 2092 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1711653199
transform 1 0 2092 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_899
timestamp 1711653199
transform 1 0 1948 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1711653199
transform 1 0 1868 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1711653199
transform 1 0 1860 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1711653199
transform 1 0 1620 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1711653199
transform 1 0 1540 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1711653199
transform 1 0 1540 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1711653199
transform 1 0 1492 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1711653199
transform 1 0 1484 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1711653199
transform 1 0 788 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1711653199
transform 1 0 708 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_909
timestamp 1711653199
transform 1 0 2908 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1711653199
transform 1 0 2556 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_911
timestamp 1711653199
transform 1 0 2516 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_912
timestamp 1711653199
transform 1 0 2468 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_913
timestamp 1711653199
transform 1 0 2292 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1711653199
transform 1 0 1924 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1711653199
transform 1 0 2972 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1711653199
transform 1 0 2868 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_917
timestamp 1711653199
transform 1 0 2868 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1711653199
transform 1 0 2324 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1711653199
transform 1 0 1596 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1711653199
transform 1 0 1596 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1711653199
transform 1 0 1388 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1711653199
transform 1 0 1380 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_923
timestamp 1711653199
transform 1 0 1300 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_924
timestamp 1711653199
transform 1 0 1204 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1711653199
transform 1 0 1164 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1711653199
transform 1 0 1100 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1711653199
transform 1 0 1060 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1711653199
transform 1 0 1028 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1711653199
transform 1 0 988 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_930
timestamp 1711653199
transform 1 0 988 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1711653199
transform 1 0 980 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1711653199
transform 1 0 980 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1711653199
transform 1 0 972 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1711653199
transform 1 0 964 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1711653199
transform 1 0 964 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1711653199
transform 1 0 948 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1711653199
transform 1 0 2564 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1711653199
transform 1 0 2508 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1711653199
transform 1 0 2444 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1711653199
transform 1 0 2876 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1711653199
transform 1 0 2788 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1711653199
transform 1 0 2676 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1711653199
transform 1 0 2396 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1711653199
transform 1 0 2372 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1711653199
transform 1 0 1860 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1711653199
transform 1 0 1676 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1711653199
transform 1 0 1676 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_948
timestamp 1711653199
transform 1 0 1660 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1711653199
transform 1 0 1652 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_950
timestamp 1711653199
transform 1 0 884 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_951
timestamp 1711653199
transform 1 0 2332 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_952
timestamp 1711653199
transform 1 0 2276 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_953
timestamp 1711653199
transform 1 0 1932 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1711653199
transform 1 0 3060 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1711653199
transform 1 0 3044 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1711653199
transform 1 0 3044 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1711653199
transform 1 0 2444 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1711653199
transform 1 0 2100 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1711653199
transform 1 0 2100 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1711653199
transform 1 0 1836 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1711653199
transform 1 0 1012 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1711653199
transform 1 0 980 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1711653199
transform 1 0 964 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_964
timestamp 1711653199
transform 1 0 964 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1711653199
transform 1 0 948 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1711653199
transform 1 0 948 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1711653199
transform 1 0 908 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1711653199
transform 1 0 892 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1711653199
transform 1 0 764 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1711653199
transform 1 0 764 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1711653199
transform 1 0 716 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1711653199
transform 1 0 716 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1711653199
transform 1 0 628 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1711653199
transform 1 0 2140 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1711653199
transform 1 0 2100 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1711653199
transform 1 0 2436 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1711653199
transform 1 0 2420 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_978
timestamp 1711653199
transform 1 0 2420 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_979
timestamp 1711653199
transform 1 0 2388 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1711653199
transform 1 0 2388 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1711653199
transform 1 0 2364 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1711653199
transform 1 0 2364 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1711653199
transform 1 0 2340 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1711653199
transform 1 0 2332 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1711653199
transform 1 0 2316 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1711653199
transform 1 0 1652 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1711653199
transform 1 0 1556 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1711653199
transform 1 0 1540 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1711653199
transform 1 0 1476 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1711653199
transform 1 0 1356 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1711653199
transform 1 0 1356 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1711653199
transform 1 0 1252 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1711653199
transform 1 0 1196 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1711653199
transform 1 0 980 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1711653199
transform 1 0 892 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1711653199
transform 1 0 884 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1711653199
transform 1 0 884 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_998
timestamp 1711653199
transform 1 0 884 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_999
timestamp 1711653199
transform 1 0 884 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1711653199
transform 1 0 884 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1711653199
transform 1 0 868 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1711653199
transform 1 0 852 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1711653199
transform 1 0 796 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1711653199
transform 1 0 692 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1711653199
transform 1 0 612 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1711653199
transform 1 0 2140 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1711653199
transform 1 0 2100 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1711653199
transform 1 0 2100 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1711653199
transform 1 0 2076 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1711653199
transform 1 0 1988 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1711653199
transform 1 0 1988 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1711653199
transform 1 0 1860 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1711653199
transform 1 0 1708 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1711653199
transform 1 0 1660 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1711653199
transform 1 0 1660 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1711653199
transform 1 0 1644 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1711653199
transform 1 0 1556 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1711653199
transform 1 0 1548 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1711653199
transform 1 0 1516 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1711653199
transform 1 0 1508 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1711653199
transform 1 0 1340 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1711653199
transform 1 0 1292 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1711653199
transform 1 0 1260 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1711653199
transform 1 0 2300 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1711653199
transform 1 0 2196 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1711653199
transform 1 0 2172 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1711653199
transform 1 0 2100 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1711653199
transform 1 0 1716 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1711653199
transform 1 0 1708 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1030
timestamp 1711653199
transform 1 0 1636 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1711653199
transform 1 0 1532 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1711653199
transform 1 0 1252 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1033
timestamp 1711653199
transform 1 0 1220 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1711653199
transform 1 0 1180 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1711653199
transform 1 0 1132 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1711653199
transform 1 0 1132 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1711653199
transform 1 0 1076 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1711653199
transform 1 0 1076 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1039
timestamp 1711653199
transform 1 0 1068 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1711653199
transform 1 0 1060 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1041
timestamp 1711653199
transform 1 0 940 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1711653199
transform 1 0 916 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_1043
timestamp 1711653199
transform 1 0 868 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_1044
timestamp 1711653199
transform 1 0 2396 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1711653199
transform 1 0 2364 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1046
timestamp 1711653199
transform 1 0 2268 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_1047
timestamp 1711653199
transform 1 0 2436 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1711653199
transform 1 0 2340 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1711653199
transform 1 0 2236 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1050
timestamp 1711653199
transform 1 0 1916 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1711653199
transform 1 0 1900 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1711653199
transform 1 0 1860 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1053
timestamp 1711653199
transform 1 0 1860 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1711653199
transform 1 0 1028 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1055
timestamp 1711653199
transform 1 0 1028 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1711653199
transform 1 0 916 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1711653199
transform 1 0 876 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1711653199
transform 1 0 812 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1711653199
transform 1 0 788 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1060
timestamp 1711653199
transform 1 0 500 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1061
timestamp 1711653199
transform 1 0 3068 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1711653199
transform 1 0 2340 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1711653199
transform 1 0 1540 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1711653199
transform 1 0 1492 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1711653199
transform 1 0 1492 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1711653199
transform 1 0 1364 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1711653199
transform 1 0 1188 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1711653199
transform 1 0 700 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1069
timestamp 1711653199
transform 1 0 508 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_1070
timestamp 1711653199
transform 1 0 500 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1071
timestamp 1711653199
transform 1 0 444 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1711653199
transform 1 0 444 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1073
timestamp 1711653199
transform 1 0 404 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1711653199
transform 1 0 380 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1711653199
transform 1 0 3292 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1711653199
transform 1 0 3260 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1711653199
transform 1 0 3260 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1711653199
transform 1 0 3228 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1079
timestamp 1711653199
transform 1 0 3228 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1080
timestamp 1711653199
transform 1 0 3204 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1711653199
transform 1 0 3148 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1711653199
transform 1 0 3148 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1083
timestamp 1711653199
transform 1 0 3084 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1084
timestamp 1711653199
transform 1 0 3084 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1711653199
transform 1 0 2972 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_1086
timestamp 1711653199
transform 1 0 2916 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1711653199
transform 1 0 2908 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1711653199
transform 1 0 2708 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1711653199
transform 1 0 2636 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1711653199
transform 1 0 2620 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1091
timestamp 1711653199
transform 1 0 1772 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1092
timestamp 1711653199
transform 1 0 1748 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1093
timestamp 1711653199
transform 1 0 1252 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1711653199
transform 1 0 1188 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1711653199
transform 1 0 1188 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1096
timestamp 1711653199
transform 1 0 1124 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1097
timestamp 1711653199
transform 1 0 588 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1711653199
transform 1 0 292 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1099
timestamp 1711653199
transform 1 0 204 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1100
timestamp 1711653199
transform 1 0 164 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_1101
timestamp 1711653199
transform 1 0 476 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1711653199
transform 1 0 420 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1711653199
transform 1 0 340 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1711653199
transform 1 0 3396 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1105
timestamp 1711653199
transform 1 0 3332 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1711653199
transform 1 0 3212 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1107
timestamp 1711653199
transform 1 0 3196 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1108
timestamp 1711653199
transform 1 0 3060 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1711653199
transform 1 0 3060 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1711653199
transform 1 0 2732 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1711653199
transform 1 0 2732 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_1112
timestamp 1711653199
transform 1 0 2508 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1711653199
transform 1 0 2516 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1711653199
transform 1 0 2404 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1711653199
transform 1 0 1132 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1711653199
transform 1 0 1036 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1117
timestamp 1711653199
transform 1 0 988 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1118
timestamp 1711653199
transform 1 0 508 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1711653199
transform 1 0 1332 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1711653199
transform 1 0 1260 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1711653199
transform 1 0 2396 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1711653199
transform 1 0 2172 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1123
timestamp 1711653199
transform 1 0 2084 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1711653199
transform 1 0 2764 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1125
timestamp 1711653199
transform 1 0 2628 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1711653199
transform 1 0 2628 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1711653199
transform 1 0 2532 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1711653199
transform 1 0 1884 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1711653199
transform 1 0 1868 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1711653199
transform 1 0 1836 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1131
timestamp 1711653199
transform 1 0 1820 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1132
timestamp 1711653199
transform 1 0 1820 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1711653199
transform 1 0 1796 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1711653199
transform 1 0 1756 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1135
timestamp 1711653199
transform 1 0 2300 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1136
timestamp 1711653199
transform 1 0 2260 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1711653199
transform 1 0 2236 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1711653199
transform 1 0 684 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1139
timestamp 1711653199
transform 1 0 652 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1711653199
transform 1 0 652 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1141
timestamp 1711653199
transform 1 0 572 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1711653199
transform 1 0 364 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1143
timestamp 1711653199
transform 1 0 740 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1711653199
transform 1 0 740 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1711653199
transform 1 0 676 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1711653199
transform 1 0 540 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1147
timestamp 1711653199
transform 1 0 3276 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1711653199
transform 1 0 3228 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1149
timestamp 1711653199
transform 1 0 3228 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1150
timestamp 1711653199
transform 1 0 3012 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_1151
timestamp 1711653199
transform 1 0 1780 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1711653199
transform 1 0 1732 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1711653199
transform 1 0 1692 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_1154
timestamp 1711653199
transform 1 0 1796 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1155
timestamp 1711653199
transform 1 0 1764 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_1156
timestamp 1711653199
transform 1 0 644 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1711653199
transform 1 0 644 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1158
timestamp 1711653199
transform 1 0 596 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1159
timestamp 1711653199
transform 1 0 596 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1160
timestamp 1711653199
transform 1 0 580 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1711653199
transform 1 0 580 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1711653199
transform 1 0 892 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1711653199
transform 1 0 812 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1164
timestamp 1711653199
transform 1 0 764 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_1165
timestamp 1711653199
transform 1 0 748 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_1166
timestamp 1711653199
transform 1 0 2540 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1167
timestamp 1711653199
transform 1 0 2260 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1711653199
transform 1 0 2260 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_1169
timestamp 1711653199
transform 1 0 1964 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1711653199
transform 1 0 3172 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1711653199
transform 1 0 3100 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1711653199
transform 1 0 3092 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1711653199
transform 1 0 3004 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1711653199
transform 1 0 3004 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1175
timestamp 1711653199
transform 1 0 3004 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_1176
timestamp 1711653199
transform 1 0 2996 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1711653199
transform 1 0 2988 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1711653199
transform 1 0 2988 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1711653199
transform 1 0 2956 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1180
timestamp 1711653199
transform 1 0 2956 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1711653199
transform 1 0 2932 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1711653199
transform 1 0 2932 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1183
timestamp 1711653199
transform 1 0 2660 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1711653199
transform 1 0 1892 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1185
timestamp 1711653199
transform 1 0 1700 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1186
timestamp 1711653199
transform 1 0 2116 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1187
timestamp 1711653199
transform 1 0 1956 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1711653199
transform 1 0 892 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1711653199
transform 1 0 796 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1190
timestamp 1711653199
transform 1 0 372 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1711653199
transform 1 0 356 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1711653199
transform 1 0 164 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1711653199
transform 1 0 1604 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1194
timestamp 1711653199
transform 1 0 1532 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1711653199
transform 1 0 1508 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1711653199
transform 1 0 1124 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1711653199
transform 1 0 332 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_1198
timestamp 1711653199
transform 1 0 324 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1199
timestamp 1711653199
transform 1 0 268 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_1200
timestamp 1711653199
transform 1 0 3348 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1201
timestamp 1711653199
transform 1 0 3300 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1711653199
transform 1 0 3284 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1711653199
transform 1 0 3108 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1711653199
transform 1 0 2932 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1205
timestamp 1711653199
transform 1 0 2908 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1711653199
transform 1 0 1892 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1207
timestamp 1711653199
transform 1 0 1860 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_1208
timestamp 1711653199
transform 1 0 1020 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1209
timestamp 1711653199
transform 1 0 804 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1711653199
transform 1 0 524 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1711653199
transform 1 0 156 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1711653199
transform 1 0 1316 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1711653199
transform 1 0 1220 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1711653199
transform 1 0 636 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1711653199
transform 1 0 588 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1711653199
transform 1 0 332 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1711653199
transform 1 0 332 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1218
timestamp 1711653199
transform 1 0 276 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1711653199
transform 1 0 3396 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1711653199
transform 1 0 3308 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1711653199
transform 1 0 3308 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1711653199
transform 1 0 2852 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1711653199
transform 1 0 2844 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1711653199
transform 1 0 2780 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1711653199
transform 1 0 2476 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1711653199
transform 1 0 2180 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1711653199
transform 1 0 2004 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1711653199
transform 1 0 1844 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1711653199
transform 1 0 1820 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1711653199
transform 1 0 1756 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1711653199
transform 1 0 1788 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1711653199
transform 1 0 1620 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1711653199
transform 1 0 1572 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1711653199
transform 1 0 1508 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1711653199
transform 1 0 1396 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1711653199
transform 1 0 404 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1711653199
transform 1 0 260 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1711653199
transform 1 0 476 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1711653199
transform 1 0 412 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_1240
timestamp 1711653199
transform 1 0 908 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1711653199
transform 1 0 804 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1711653199
transform 1 0 2308 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1243
timestamp 1711653199
transform 1 0 2276 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1711653199
transform 1 0 2220 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1245
timestamp 1711653199
transform 1 0 2492 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1711653199
transform 1 0 2324 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1711653199
transform 1 0 2428 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1248
timestamp 1711653199
transform 1 0 2388 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1711653199
transform 1 0 2684 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1711653199
transform 1 0 2452 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1251
timestamp 1711653199
transform 1 0 3284 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1711653199
transform 1 0 3140 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1711653199
transform 1 0 3108 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1711653199
transform 1 0 3356 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1711653199
transform 1 0 3252 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1711653199
transform 1 0 3132 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1711653199
transform 1 0 3364 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1711653199
transform 1 0 3252 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1711653199
transform 1 0 3364 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1711653199
transform 1 0 3332 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1711653199
transform 1 0 3228 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1711653199
transform 1 0 3140 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1711653199
transform 1 0 2980 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1711653199
transform 1 0 2924 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1711653199
transform 1 0 2876 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1711653199
transform 1 0 3236 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1711653199
transform 1 0 3204 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1711653199
transform 1 0 3180 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1711653199
transform 1 0 3252 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1711653199
transform 1 0 3220 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1271
timestamp 1711653199
transform 1 0 3188 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1711653199
transform 1 0 3028 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1711653199
transform 1 0 2980 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1711653199
transform 1 0 2404 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1711653199
transform 1 0 2380 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1711653199
transform 1 0 2196 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1277
timestamp 1711653199
transform 1 0 3228 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1711653199
transform 1 0 3084 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1711653199
transform 1 0 1140 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1711653199
transform 1 0 1084 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1711653199
transform 1 0 1084 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1711653199
transform 1 0 1068 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1711653199
transform 1 0 2412 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1711653199
transform 1 0 2324 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1711653199
transform 1 0 3036 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1286
timestamp 1711653199
transform 1 0 2932 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1711653199
transform 1 0 3364 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1711653199
transform 1 0 3324 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1711653199
transform 1 0 3356 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1290
timestamp 1711653199
transform 1 0 3332 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1711653199
transform 1 0 3340 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1711653199
transform 1 0 3116 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_1293
timestamp 1711653199
transform 1 0 3396 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1711653199
transform 1 0 3324 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1711653199
transform 1 0 3244 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1296
timestamp 1711653199
transform 1 0 3196 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1711653199
transform 1 0 3172 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1711653199
transform 1 0 1420 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1711653199
transform 1 0 1372 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_1300
timestamp 1711653199
transform 1 0 2756 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1711653199
transform 1 0 2692 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1711653199
transform 1 0 2668 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_1303
timestamp 1711653199
transform 1 0 2724 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1711653199
transform 1 0 2676 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1711653199
transform 1 0 2012 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1711653199
transform 1 0 2100 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1711653199
transform 1 0 1956 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_1308
timestamp 1711653199
transform 1 0 1444 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1711653199
transform 1 0 1740 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1711653199
transform 1 0 1492 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1711653199
transform 1 0 2332 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1711653199
transform 1 0 2308 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1711653199
transform 1 0 2308 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1314
timestamp 1711653199
transform 1 0 2300 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1711653199
transform 1 0 2212 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1711653199
transform 1 0 2212 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1711653199
transform 1 0 2204 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1711653199
transform 1 0 2060 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1711653199
transform 1 0 2516 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1711653199
transform 1 0 2468 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1711653199
transform 1 0 2372 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1322
timestamp 1711653199
transform 1 0 2340 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1711653199
transform 1 0 2364 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1711653199
transform 1 0 2284 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1711653199
transform 1 0 2244 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_1326
timestamp 1711653199
transform 1 0 2604 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1327
timestamp 1711653199
transform 1 0 2564 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1328
timestamp 1711653199
transform 1 0 2284 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1711653199
transform 1 0 2012 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1711653199
transform 1 0 1980 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1711653199
transform 1 0 2364 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1332
timestamp 1711653199
transform 1 0 2324 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_1333
timestamp 1711653199
transform 1 0 2532 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1711653199
transform 1 0 2380 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1711653199
transform 1 0 2564 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1336
timestamp 1711653199
transform 1 0 2148 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_1337
timestamp 1711653199
transform 1 0 2140 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1338
timestamp 1711653199
transform 1 0 2076 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1711653199
transform 1 0 2148 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1340
timestamp 1711653199
transform 1 0 2084 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_1341
timestamp 1711653199
transform 1 0 2508 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1711653199
transform 1 0 1932 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1711653199
transform 1 0 1684 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1711653199
transform 1 0 1532 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1345
timestamp 1711653199
transform 1 0 1532 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1711653199
transform 1 0 1292 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1711653199
transform 1 0 2228 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1711653199
transform 1 0 1820 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1349
timestamp 1711653199
transform 1 0 1820 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1711653199
transform 1 0 1796 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1351
timestamp 1711653199
transform 1 0 1148 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1711653199
transform 1 0 1052 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1353
timestamp 1711653199
transform 1 0 756 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1711653199
transform 1 0 684 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_1355
timestamp 1711653199
transform 1 0 644 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1711653199
transform 1 0 604 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1357
timestamp 1711653199
transform 1 0 772 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1711653199
transform 1 0 700 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_1359
timestamp 1711653199
transform 1 0 252 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1711653199
transform 1 0 228 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1711653199
transform 1 0 332 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1711653199
transform 1 0 260 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1711653199
transform 1 0 260 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1711653199
transform 1 0 228 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1711653199
transform 1 0 196 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1711653199
transform 1 0 164 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1711653199
transform 1 0 116 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1711653199
transform 1 0 180 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1711653199
transform 1 0 132 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1711653199
transform 1 0 132 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1711653199
transform 1 0 132 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1711653199
transform 1 0 100 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1711653199
transform 1 0 100 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1374
timestamp 1711653199
transform 1 0 92 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_1375
timestamp 1711653199
transform 1 0 860 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1711653199
transform 1 0 708 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1711653199
transform 1 0 676 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1711653199
transform 1 0 644 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1711653199
transform 1 0 996 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1711653199
transform 1 0 948 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1711653199
transform 1 0 916 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1382
timestamp 1711653199
transform 1 0 1260 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1711653199
transform 1 0 1220 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1711653199
transform 1 0 972 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1711653199
transform 1 0 948 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1711653199
transform 1 0 892 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1711653199
transform 1 0 828 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1388
timestamp 1711653199
transform 1 0 828 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_1389
timestamp 1711653199
transform 1 0 708 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1711653199
transform 1 0 852 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1391
timestamp 1711653199
transform 1 0 812 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1711653199
transform 1 0 652 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1711653199
transform 1 0 596 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1711653199
transform 1 0 1252 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1711653199
transform 1 0 644 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1711653199
transform 1 0 580 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1711653199
transform 1 0 580 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_1398
timestamp 1711653199
transform 1 0 492 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1399
timestamp 1711653199
transform 1 0 444 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1711653199
transform 1 0 1116 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1711653199
transform 1 0 876 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1711653199
transform 1 0 860 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_1403
timestamp 1711653199
transform 1 0 596 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1711653199
transform 1 0 996 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1711653199
transform 1 0 756 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1711653199
transform 1 0 1092 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1711653199
transform 1 0 956 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1711653199
transform 1 0 1052 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1711653199
transform 1 0 996 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1711653199
transform 1 0 1052 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1711653199
transform 1 0 908 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1711653199
transform 1 0 964 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1711653199
transform 1 0 892 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1414
timestamp 1711653199
transform 1 0 892 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1711653199
transform 1 0 772 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1711653199
transform 1 0 428 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1711653199
transform 1 0 364 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_1418
timestamp 1711653199
transform 1 0 124 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1711653199
transform 1 0 76 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_1420
timestamp 1711653199
transform 1 0 228 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_1421
timestamp 1711653199
transform 1 0 164 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1422
timestamp 1711653199
transform 1 0 132 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_1423
timestamp 1711653199
transform 1 0 1124 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1424
timestamp 1711653199
transform 1 0 1060 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1711653199
transform 1 0 1116 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1426
timestamp 1711653199
transform 1 0 1068 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1711653199
transform 1 0 1876 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1428
timestamp 1711653199
transform 1 0 1804 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1429
timestamp 1711653199
transform 1 0 1756 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1711653199
transform 1 0 1692 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1431
timestamp 1711653199
transform 1 0 1556 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1711653199
transform 1 0 1428 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1433
timestamp 1711653199
transform 1 0 1140 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1434
timestamp 1711653199
transform 1 0 1900 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1711653199
transform 1 0 1860 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1436
timestamp 1711653199
transform 1 0 1796 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1711653199
transform 1 0 1580 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1711653199
transform 1 0 2284 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1711653199
transform 1 0 2236 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1711653199
transform 1 0 2124 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1441
timestamp 1711653199
transform 1 0 2420 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1711653199
transform 1 0 2276 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1711653199
transform 1 0 2276 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1444
timestamp 1711653199
transform 1 0 2156 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1711653199
transform 1 0 2116 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1711653199
transform 1 0 1988 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1711653199
transform 1 0 1660 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1711653199
transform 1 0 1444 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1711653199
transform 1 0 3028 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1711653199
transform 1 0 2972 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1711653199
transform 1 0 2940 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1711653199
transform 1 0 3364 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_1453
timestamp 1711653199
transform 1 0 3364 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1711653199
transform 1 0 3308 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_1455
timestamp 1711653199
transform 1 0 3284 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1711653199
transform 1 0 3252 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1711653199
transform 1 0 3380 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1711653199
transform 1 0 3308 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1711653199
transform 1 0 3380 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1711653199
transform 1 0 3356 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1711653199
transform 1 0 3268 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1462
timestamp 1711653199
transform 1 0 3380 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1711653199
transform 1 0 3300 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1711653199
transform 1 0 2948 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1711653199
transform 1 0 2868 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1711653199
transform 1 0 2492 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1711653199
transform 1 0 2396 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1711653199
transform 1 0 2364 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1711653199
transform 1 0 2324 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1711653199
transform 1 0 2620 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1471
timestamp 1711653199
transform 1 0 2548 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1711653199
transform 1 0 2444 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1711653199
transform 1 0 2364 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1711653199
transform 1 0 2292 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1711653199
transform 1 0 2276 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1476
timestamp 1711653199
transform 1 0 2220 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_1477
timestamp 1711653199
transform 1 0 2756 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1711653199
transform 1 0 2724 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_1479
timestamp 1711653199
transform 1 0 2972 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1480
timestamp 1711653199
transform 1 0 2828 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1481
timestamp 1711653199
transform 1 0 1892 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1711653199
transform 1 0 1764 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1711653199
transform 1 0 1660 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1484
timestamp 1711653199
transform 1 0 1532 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1485
timestamp 1711653199
transform 1 0 1396 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1711653199
transform 1 0 1292 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1487
timestamp 1711653199
transform 1 0 1156 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1488
timestamp 1711653199
transform 1 0 1020 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1711653199
transform 1 0 876 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1711653199
transform 1 0 580 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1711653199
transform 1 0 468 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1711653199
transform 1 0 316 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1711653199
transform 1 0 3204 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1711653199
transform 1 0 2836 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1711653199
transform 1 0 2820 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1711653199
transform 1 0 2732 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1711653199
transform 1 0 2628 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1711653199
transform 1 0 2612 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1711653199
transform 1 0 1884 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1711653199
transform 1 0 1884 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1711653199
transform 1 0 1716 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1711653199
transform 1 0 1716 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1711653199
transform 1 0 1564 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1711653199
transform 1 0 1556 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1711653199
transform 1 0 1500 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1711653199
transform 1 0 1500 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1507
timestamp 1711653199
transform 1 0 1460 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_1508
timestamp 1711653199
transform 1 0 1452 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_1509
timestamp 1711653199
transform 1 0 1268 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1510
timestamp 1711653199
transform 1 0 788 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1711653199
transform 1 0 564 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1512
timestamp 1711653199
transform 1 0 564 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1513
timestamp 1711653199
transform 1 0 420 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1711653199
transform 1 0 420 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1711653199
transform 1 0 308 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1711653199
transform 1 0 276 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1517
timestamp 1711653199
transform 1 0 276 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1518
timestamp 1711653199
transform 1 0 172 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_1519
timestamp 1711653199
transform 1 0 92 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1520
timestamp 1711653199
transform 1 0 3316 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1521
timestamp 1711653199
transform 1 0 3316 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1711653199
transform 1 0 3268 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1711653199
transform 1 0 3268 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1524
timestamp 1711653199
transform 1 0 3220 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1711653199
transform 1 0 3004 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1526
timestamp 1711653199
transform 1 0 3004 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1711653199
transform 1 0 2812 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1528
timestamp 1711653199
transform 1 0 2748 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_1529
timestamp 1711653199
transform 1 0 2732 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1530
timestamp 1711653199
transform 1 0 2644 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_1531
timestamp 1711653199
transform 1 0 2644 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1711653199
transform 1 0 2596 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1533
timestamp 1711653199
transform 1 0 2564 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1534
timestamp 1711653199
transform 1 0 2468 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1711653199
transform 1 0 3308 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1711653199
transform 1 0 3092 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1537
timestamp 1711653199
transform 1 0 2900 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1711653199
transform 1 0 2900 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1711653199
transform 1 0 2804 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1540
timestamp 1711653199
transform 1 0 2788 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1541
timestamp 1711653199
transform 1 0 2716 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1711653199
transform 1 0 2508 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1711653199
transform 1 0 2372 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1711653199
transform 1 0 2276 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1711653199
transform 1 0 2172 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1711653199
transform 1 0 2076 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1711653199
transform 1 0 1972 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1711653199
transform 1 0 1972 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1711653199
transform 1 0 1900 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1550
timestamp 1711653199
transform 1 0 1924 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1711653199
transform 1 0 1844 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1711653199
transform 1 0 1812 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1711653199
transform 1 0 1812 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1711653199
transform 1 0 1708 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1711653199
transform 1 0 1708 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1556
timestamp 1711653199
transform 1 0 1572 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1711653199
transform 1 0 1468 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1711653199
transform 1 0 1300 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1711653199
transform 1 0 1004 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1711653199
transform 1 0 1004 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1711653199
transform 1 0 916 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1711653199
transform 1 0 916 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1711653199
transform 1 0 820 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1711653199
transform 1 0 692 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1711653199
transform 1 0 580 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1711653199
transform 1 0 428 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1567
timestamp 1711653199
transform 1 0 428 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1711653199
transform 1 0 380 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1711653199
transform 1 0 276 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1711653199
transform 1 0 1964 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1711653199
transform 1 0 1860 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1711653199
transform 1 0 1860 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1573
timestamp 1711653199
transform 1 0 1828 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1574
timestamp 1711653199
transform 1 0 1828 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1711653199
transform 1 0 1780 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1711653199
transform 1 0 1724 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1711653199
transform 1 0 1508 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1711653199
transform 1 0 980 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_1579
timestamp 1711653199
transform 1 0 980 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1711653199
transform 1 0 732 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1711653199
transform 1 0 420 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1711653199
transform 1 0 340 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1711653199
transform 1 0 340 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1711653199
transform 1 0 204 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1711653199
transform 1 0 156 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1711653199
transform 1 0 156 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1587
timestamp 1711653199
transform 1 0 92 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1711653199
transform 1 0 92 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1711653199
transform 1 0 2556 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1711653199
transform 1 0 2444 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1711653199
transform 1 0 2340 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1711653199
transform 1 0 2300 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1711653199
transform 1 0 2236 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1711653199
transform 1 0 2196 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1711653199
transform 1 0 2196 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1711653199
transform 1 0 2036 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1711653199
transform 1 0 1628 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1711653199
transform 1 0 1516 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1711653199
transform 1 0 1476 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1711653199
transform 1 0 1412 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1711653199
transform 1 0 1364 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1711653199
transform 1 0 1244 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1711653199
transform 1 0 1156 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1604
timestamp 1711653199
transform 1 0 1044 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1711653199
transform 1 0 844 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1606
timestamp 1711653199
transform 1 0 812 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1711653199
transform 1 0 692 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1711653199
transform 1 0 572 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1711653199
transform 1 0 524 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1610
timestamp 1711653199
transform 1 0 460 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1711653199
transform 1 0 412 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1711653199
transform 1 0 308 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1711653199
transform 1 0 196 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1711653199
transform 1 0 92 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1711653199
transform 1 0 3180 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1711653199
transform 1 0 3164 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1711653199
transform 1 0 3068 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1711653199
transform 1 0 2980 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1711653199
transform 1 0 2916 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1711653199
transform 1 0 2908 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1711653199
transform 1 0 2876 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1711653199
transform 1 0 2868 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1711653199
transform 1 0 2844 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1711653199
transform 1 0 2140 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1711653199
transform 1 0 2140 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1711653199
transform 1 0 2036 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1711653199
transform 1 0 1932 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1711653199
transform 1 0 1932 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1711653199
transform 1 0 1788 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1711653199
transform 1 0 1788 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1711653199
transform 1 0 1516 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1711653199
transform 1 0 1476 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1711653199
transform 1 0 1356 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1711653199
transform 1 0 1860 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1711653199
transform 1 0 1812 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1636
timestamp 1711653199
transform 1 0 1780 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1711653199
transform 1 0 1476 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1638
timestamp 1711653199
transform 1 0 1460 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1639
timestamp 1711653199
transform 1 0 1228 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1711653199
transform 1 0 2612 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1711653199
transform 1 0 2588 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1642
timestamp 1711653199
transform 1 0 2484 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1643
timestamp 1711653199
transform 1 0 3284 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1711653199
transform 1 0 3060 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1711653199
transform 1 0 2924 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1646
timestamp 1711653199
transform 1 0 2620 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1711653199
transform 1 0 2596 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1711653199
transform 1 0 2764 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1711653199
transform 1 0 2660 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1711653199
transform 1 0 2612 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_1651
timestamp 1711653199
transform 1 0 2604 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1652
timestamp 1711653199
transform 1 0 2604 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1653
timestamp 1711653199
transform 1 0 2572 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_1654
timestamp 1711653199
transform 1 0 2572 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1711653199
transform 1 0 2524 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1711653199
transform 1 0 2460 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1711653199
transform 1 0 3276 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_1658
timestamp 1711653199
transform 1 0 3052 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1711653199
transform 1 0 3012 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1711653199
transform 1 0 2988 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1661
timestamp 1711653199
transform 1 0 2988 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1662
timestamp 1711653199
transform 1 0 2940 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_1663
timestamp 1711653199
transform 1 0 2860 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1711653199
transform 1 0 2860 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_1665
timestamp 1711653199
transform 1 0 2852 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_1666
timestamp 1711653199
transform 1 0 2852 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_1667
timestamp 1711653199
transform 1 0 2740 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1711653199
transform 1 0 2564 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1711653199
transform 1 0 2028 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1711653199
transform 1 0 2012 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1711653199
transform 1 0 1932 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_1672
timestamp 1711653199
transform 1 0 1932 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1673
timestamp 1711653199
transform 1 0 1780 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1711653199
transform 1 0 1484 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1675
timestamp 1711653199
transform 1 0 1028 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1711653199
transform 1 0 1028 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1677
timestamp 1711653199
transform 1 0 932 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1711653199
transform 1 0 668 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1711653199
transform 1 0 668 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1711653199
transform 1 0 516 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1711653199
transform 1 0 516 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1682
timestamp 1711653199
transform 1 0 364 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1711653199
transform 1 0 364 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1711653199
transform 1 0 260 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1685
timestamp 1711653199
transform 1 0 228 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1711653199
transform 1 0 212 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1687
timestamp 1711653199
transform 1 0 204 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_1688
timestamp 1711653199
transform 1 0 196 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_1689
timestamp 1711653199
transform 1 0 2124 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1711653199
transform 1 0 2028 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1711653199
transform 1 0 1908 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1692
timestamp 1711653199
transform 1 0 1836 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1711653199
transform 1 0 1740 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1694
timestamp 1711653199
transform 1 0 1948 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1711653199
transform 1 0 1852 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1696
timestamp 1711653199
transform 1 0 1668 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1711653199
transform 1 0 1636 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1698
timestamp 1711653199
transform 1 0 1756 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1699
timestamp 1711653199
transform 1 0 1388 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1711653199
transform 1 0 1388 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1701
timestamp 1711653199
transform 1 0 1324 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1702
timestamp 1711653199
transform 1 0 932 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1703
timestamp 1711653199
transform 1 0 828 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1711653199
transform 1 0 764 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1705
timestamp 1711653199
transform 1 0 572 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_1706
timestamp 1711653199
transform 1 0 2348 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1711653199
transform 1 0 1940 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1711653199
transform 1 0 1844 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_1709
timestamp 1711653199
transform 1 0 1788 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1711653199
transform 1 0 500 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_1711
timestamp 1711653199
transform 1 0 436 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1711653199
transform 1 0 404 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1711653199
transform 1 0 292 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1711653199
transform 1 0 252 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1711653199
transform 1 0 212 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1711653199
transform 1 0 204 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1711653199
transform 1 0 124 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1718
timestamp 1711653199
transform 1 0 2148 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1711653199
transform 1 0 2060 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1711653199
transform 1 0 2052 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1711653199
transform 1 0 1868 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1711653199
transform 1 0 1868 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_1723
timestamp 1711653199
transform 1 0 1612 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1711653199
transform 1 0 1260 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1711653199
transform 1 0 1156 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1711653199
transform 1 0 1156 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_1727
timestamp 1711653199
transform 1 0 1132 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1728
timestamp 1711653199
transform 1 0 1092 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_1729
timestamp 1711653199
transform 1 0 2652 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1711653199
transform 1 0 2532 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1731
timestamp 1711653199
transform 1 0 2284 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1711653199
transform 1 0 2164 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_1733
timestamp 1711653199
transform 1 0 1892 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1734
timestamp 1711653199
transform 1 0 1860 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1711653199
transform 1 0 1684 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1711653199
transform 1 0 1588 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1711653199
transform 1 0 2180 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1711653199
transform 1 0 2140 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1711653199
transform 1 0 2116 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1711653199
transform 1 0 2092 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1711653199
transform 1 0 1988 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1711653199
transform 1 0 1892 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1711653199
transform 1 0 1820 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1711653199
transform 1 0 1812 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1745
timestamp 1711653199
transform 1 0 1652 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1711653199
transform 1 0 1636 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_1747
timestamp 1711653199
transform 1 0 1428 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1748
timestamp 1711653199
transform 1 0 1364 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1711653199
transform 1 0 1300 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1711653199
transform 1 0 1244 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1711653199
transform 1 0 1244 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1711653199
transform 1 0 1212 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1711653199
transform 1 0 1204 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1711653199
transform 1 0 1148 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1711653199
transform 1 0 948 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1711653199
transform 1 0 948 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1711653199
transform 1 0 884 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1711653199
transform 1 0 884 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1711653199
transform 1 0 820 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1711653199
transform 1 0 628 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1711653199
transform 1 0 628 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1711653199
transform 1 0 372 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1763
timestamp 1711653199
transform 1 0 252 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1711653199
transform 1 0 2684 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1711653199
transform 1 0 2668 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1711653199
transform 1 0 2604 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1711653199
transform 1 0 2364 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1711653199
transform 1 0 2716 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1711653199
transform 1 0 2476 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1711653199
transform 1 0 2228 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1711653199
transform 1 0 1988 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_1772
timestamp 1711653199
transform 1 0 2348 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1711653199
transform 1 0 2332 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1711653199
transform 1 0 2308 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_1775
timestamp 1711653199
transform 1 0 2308 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_1776
timestamp 1711653199
transform 1 0 2172 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_1777
timestamp 1711653199
transform 1 0 2172 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_1778
timestamp 1711653199
transform 1 0 2092 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1711653199
transform 1 0 2092 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_1780
timestamp 1711653199
transform 1 0 1804 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1711653199
transform 1 0 1724 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1711653199
transform 1 0 1716 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1783
timestamp 1711653199
transform 1 0 1692 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_1784
timestamp 1711653199
transform 1 0 1684 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_1785
timestamp 1711653199
transform 1 0 1676 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_1786
timestamp 1711653199
transform 1 0 1676 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1787
timestamp 1711653199
transform 1 0 1652 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1711653199
transform 1 0 1556 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1711653199
transform 1 0 1556 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1711653199
transform 1 0 1460 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1711653199
transform 1 0 1372 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1711653199
transform 1 0 1220 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1793
timestamp 1711653199
transform 1 0 1100 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1711653199
transform 1 0 1020 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_1795
timestamp 1711653199
transform 1 0 940 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1796
timestamp 1711653199
transform 1 0 724 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1711653199
transform 1 0 628 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1711653199
transform 1 0 604 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1711653199
transform 1 0 604 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1711653199
transform 1 0 588 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1801
timestamp 1711653199
transform 1 0 564 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1711653199
transform 1 0 556 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1711653199
transform 1 0 524 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1804
timestamp 1711653199
transform 1 0 508 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1711653199
transform 1 0 492 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1711653199
transform 1 0 492 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1711653199
transform 1 0 468 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1711653199
transform 1 0 468 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1711653199
transform 1 0 444 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1711653199
transform 1 0 2316 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1711653199
transform 1 0 2204 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1711653199
transform 1 0 2204 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1711653199
transform 1 0 2140 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1711653199
transform 1 0 2036 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1711653199
transform 1 0 1956 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1711653199
transform 1 0 1836 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1711653199
transform 1 0 1812 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1711653199
transform 1 0 1804 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1819
timestamp 1711653199
transform 1 0 1708 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1711653199
transform 1 0 1700 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1711653199
transform 1 0 1588 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1711653199
transform 1 0 1556 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1711653199
transform 1 0 1540 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1824
timestamp 1711653199
transform 1 0 1540 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1711653199
transform 1 0 1436 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1711653199
transform 1 0 1388 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1711653199
transform 1 0 1308 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1711653199
transform 1 0 1140 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_1829
timestamp 1711653199
transform 1 0 1020 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1830
timestamp 1711653199
transform 1 0 916 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1711653199
transform 1 0 908 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1711653199
transform 1 0 900 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1833
timestamp 1711653199
transform 1 0 692 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1711653199
transform 1 0 676 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1711653199
transform 1 0 676 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1711653199
transform 1 0 532 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1711653199
transform 1 0 532 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1711653199
transform 1 0 492 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1839
timestamp 1711653199
transform 1 0 412 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1711653199
transform 1 0 364 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1711653199
transform 1 0 332 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1711653199
transform 1 0 252 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1711653199
transform 1 0 236 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1711653199
transform 1 0 3188 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1711653199
transform 1 0 3156 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1711653199
transform 1 0 3108 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1711653199
transform 1 0 3108 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1711653199
transform 1 0 3068 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1711653199
transform 1 0 3052 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1711653199
transform 1 0 2684 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_1851
timestamp 1711653199
transform 1 0 2260 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1711653199
transform 1 0 3012 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1853
timestamp 1711653199
transform 1 0 2988 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1711653199
transform 1 0 2916 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1855
timestamp 1711653199
transform 1 0 3300 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1711653199
transform 1 0 3100 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1711653199
transform 1 0 3092 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1711653199
transform 1 0 2644 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1711653199
transform 1 0 2308 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1711653199
transform 1 0 2260 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1711653199
transform 1 0 2244 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1711653199
transform 1 0 2236 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1711653199
transform 1 0 2188 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1711653199
transform 1 0 2180 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1865
timestamp 1711653199
transform 1 0 2124 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1711653199
transform 1 0 2100 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1711653199
transform 1 0 2068 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1711653199
transform 1 0 2060 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1711653199
transform 1 0 2060 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1711653199
transform 1 0 2028 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1711653199
transform 1 0 2020 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1711653199
transform 1 0 2020 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1711653199
transform 1 0 2012 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1874
timestamp 1711653199
transform 1 0 1948 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1711653199
transform 1 0 1636 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_1876
timestamp 1711653199
transform 1 0 1580 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1711653199
transform 1 0 1388 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1711653199
transform 1 0 1220 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1711653199
transform 1 0 1132 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1711653199
transform 1 0 1116 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1711653199
transform 1 0 988 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1711653199
transform 1 0 980 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1711653199
transform 1 0 948 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1711653199
transform 1 0 948 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1711653199
transform 1 0 884 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1711653199
transform 1 0 884 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1711653199
transform 1 0 844 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1711653199
transform 1 0 700 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_1889
timestamp 1711653199
transform 1 0 692 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1711653199
transform 1 0 668 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1711653199
transform 1 0 628 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1711653199
transform 1 0 628 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1711653199
transform 1 0 612 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1711653199
transform 1 0 388 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1711653199
transform 1 0 252 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1711653199
transform 1 0 236 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1711653199
transform 1 0 172 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_1898
timestamp 1711653199
transform 1 0 3028 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1711653199
transform 1 0 2988 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_1900
timestamp 1711653199
transform 1 0 2916 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1711653199
transform 1 0 2756 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1711653199
transform 1 0 2580 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1903
timestamp 1711653199
transform 1 0 2556 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1711653199
transform 1 0 2444 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1711653199
transform 1 0 2276 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1906
timestamp 1711653199
transform 1 0 2228 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1711653199
transform 1 0 2140 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1711653199
transform 1 0 3316 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1711653199
transform 1 0 3308 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1910
timestamp 1711653199
transform 1 0 3300 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1711653199
transform 1 0 3252 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1912
timestamp 1711653199
transform 1 0 3252 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1913
timestamp 1711653199
transform 1 0 3156 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1711653199
transform 1 0 3100 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1711653199
transform 1 0 3100 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1916
timestamp 1711653199
transform 1 0 3044 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1711653199
transform 1 0 3044 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1711653199
transform 1 0 3028 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1711653199
transform 1 0 3028 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1711653199
transform 1 0 2956 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1711653199
transform 1 0 2956 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1711653199
transform 1 0 2940 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_1923
timestamp 1711653199
transform 1 0 2708 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1711653199
transform 1 0 2564 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1925
timestamp 1711653199
transform 1 0 2012 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_1926
timestamp 1711653199
transform 1 0 1964 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1711653199
transform 1 0 1908 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1711653199
transform 1 0 1732 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1711653199
transform 1 0 1692 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1930
timestamp 1711653199
transform 1 0 1652 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1711653199
transform 1 0 1652 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1711653199
transform 1 0 1644 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_1933
timestamp 1711653199
transform 1 0 1604 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1711653199
transform 1 0 1524 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1711653199
transform 1 0 1492 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1711653199
transform 1 0 1428 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1711653199
transform 1 0 1284 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1711653199
transform 1 0 1284 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1711653199
transform 1 0 1036 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1940
timestamp 1711653199
transform 1 0 988 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1941
timestamp 1711653199
transform 1 0 796 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1711653199
transform 1 0 796 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1943
timestamp 1711653199
transform 1 0 748 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1711653199
transform 1 0 644 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_1945
timestamp 1711653199
transform 1 0 644 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_1946
timestamp 1711653199
transform 1 0 524 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1711653199
transform 1 0 380 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1711653199
transform 1 0 372 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1711653199
transform 1 0 324 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_1950
timestamp 1711653199
transform 1 0 244 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1711653199
transform 1 0 244 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_1952
timestamp 1711653199
transform 1 0 196 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1953
timestamp 1711653199
transform 1 0 3188 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1711653199
transform 1 0 3164 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1711653199
transform 1 0 2804 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1711653199
transform 1 0 3252 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1711653199
transform 1 0 3252 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1711653199
transform 1 0 3188 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1711653199
transform 1 0 2876 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1711653199
transform 1 0 2700 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1711653199
transform 1 0 3180 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1711653199
transform 1 0 3180 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1711653199
transform 1 0 3180 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1711653199
transform 1 0 3132 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1711653199
transform 1 0 2644 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1711653199
transform 1 0 2636 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1967
timestamp 1711653199
transform 1 0 2516 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_1968
timestamp 1711653199
transform 1 0 2516 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1969
timestamp 1711653199
transform 1 0 1700 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1711653199
transform 1 0 1628 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1711653199
transform 1 0 1628 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1711653199
transform 1 0 1348 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_1973
timestamp 1711653199
transform 1 0 1348 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1711653199
transform 1 0 1228 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1711653199
transform 1 0 1228 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1976
timestamp 1711653199
transform 1 0 996 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1711653199
transform 1 0 916 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1711653199
transform 1 0 908 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1711653199
transform 1 0 764 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1711653199
transform 1 0 764 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1981
timestamp 1711653199
transform 1 0 692 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1982
timestamp 1711653199
transform 1 0 484 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1711653199
transform 1 0 476 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1711653199
transform 1 0 348 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1711653199
transform 1 0 292 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1711653199
transform 1 0 3300 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1711653199
transform 1 0 3292 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1711653199
transform 1 0 3260 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1711653199
transform 1 0 3236 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1711653199
transform 1 0 3236 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1711653199
transform 1 0 3060 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_1992
timestamp 1711653199
transform 1 0 3060 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1711653199
transform 1 0 3060 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1711653199
transform 1 0 3028 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1711653199
transform 1 0 2956 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1711653199
transform 1 0 2372 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1997
timestamp 1711653199
transform 1 0 2276 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_1998
timestamp 1711653199
transform 1 0 2116 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1711653199
transform 1 0 1996 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1711653199
transform 1 0 1996 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1711653199
transform 1 0 1900 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2002
timestamp 1711653199
transform 1 0 1868 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1711653199
transform 1 0 1844 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1711653199
transform 1 0 1788 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1711653199
transform 1 0 1788 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1711653199
transform 1 0 1620 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1711653199
transform 1 0 1620 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1711653199
transform 1 0 1580 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1711653199
transform 1 0 1572 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1711653199
transform 1 0 604 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1711653199
transform 1 0 516 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1711653199
transform 1 0 516 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1711653199
transform 1 0 444 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1711653199
transform 1 0 444 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1711653199
transform 1 0 332 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1711653199
transform 1 0 204 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1711653199
transform 1 0 196 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2018
timestamp 1711653199
transform 1 0 164 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2019
timestamp 1711653199
transform 1 0 3132 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1711653199
transform 1 0 3108 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_2021
timestamp 1711653199
transform 1 0 3116 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1711653199
transform 1 0 2492 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1711653199
transform 1 0 2396 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1711653199
transform 1 0 3260 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1711653199
transform 1 0 3260 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1711653199
transform 1 0 3220 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2027
timestamp 1711653199
transform 1 0 3220 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1711653199
transform 1 0 3140 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2029
timestamp 1711653199
transform 1 0 3140 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1711653199
transform 1 0 3140 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2031
timestamp 1711653199
transform 1 0 3116 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1711653199
transform 1 0 3108 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1711653199
transform 1 0 3028 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2034
timestamp 1711653199
transform 1 0 2972 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_2035
timestamp 1711653199
transform 1 0 2956 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2036
timestamp 1711653199
transform 1 0 2748 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2037
timestamp 1711653199
transform 1 0 2748 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2038
timestamp 1711653199
transform 1 0 2508 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1711653199
transform 1 0 2460 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2040
timestamp 1711653199
transform 1 0 2292 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1711653199
transform 1 0 2204 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_2042
timestamp 1711653199
transform 1 0 1996 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1711653199
transform 1 0 1996 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2044
timestamp 1711653199
transform 1 0 1924 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1711653199
transform 1 0 1788 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2046
timestamp 1711653199
transform 1 0 1788 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1711653199
transform 1 0 1484 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2048
timestamp 1711653199
transform 1 0 1484 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1711653199
transform 1 0 1484 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1711653199
transform 1 0 1348 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2051
timestamp 1711653199
transform 1 0 1316 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1711653199
transform 1 0 1116 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1711653199
transform 1 0 1100 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2054
timestamp 1711653199
transform 1 0 1100 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2055
timestamp 1711653199
transform 1 0 908 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1711653199
transform 1 0 892 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1711653199
transform 1 0 780 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1711653199
transform 1 0 780 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1711653199
transform 1 0 588 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1711653199
transform 1 0 588 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1711653199
transform 1 0 484 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1711653199
transform 1 0 436 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1711653199
transform 1 0 436 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1711653199
transform 1 0 332 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1711653199
transform 1 0 180 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2066
timestamp 1711653199
transform 1 0 172 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2067
timestamp 1711653199
transform 1 0 140 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1711653199
transform 1 0 140 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1711653199
transform 1 0 2628 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2070
timestamp 1711653199
transform 1 0 2380 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1711653199
transform 1 0 2252 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1711653199
transform 1 0 2100 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1711653199
transform 1 0 2100 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1711653199
transform 1 0 1956 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2075
timestamp 1711653199
transform 1 0 1940 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1711653199
transform 1 0 1876 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2077
timestamp 1711653199
transform 1 0 1724 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2078
timestamp 1711653199
transform 1 0 1508 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2079
timestamp 1711653199
transform 1 0 1508 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1711653199
transform 1 0 1244 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1711653199
transform 1 0 1052 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1711653199
transform 1 0 1020 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1711653199
transform 1 0 1020 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1711653199
transform 1 0 548 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2085
timestamp 1711653199
transform 1 0 420 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1711653199
transform 1 0 420 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1711653199
transform 1 0 404 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1711653199
transform 1 0 404 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1711653199
transform 1 0 3316 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1711653199
transform 1 0 3124 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1711653199
transform 1 0 2796 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1711653199
transform 1 0 2356 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1711653199
transform 1 0 2348 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1711653199
transform 1 0 1356 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1711653199
transform 1 0 924 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1711653199
transform 1 0 628 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1711653199
transform 1 0 420 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1711653199
transform 1 0 372 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1711653199
transform 1 0 260 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1711653199
transform 1 0 244 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1711653199
transform 1 0 172 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1711653199
transform 1 0 140 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1711653199
transform 1 0 2972 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1711653199
transform 1 0 2876 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1711653199
transform 1 0 3156 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1711653199
transform 1 0 3124 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1711653199
transform 1 0 2940 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1711653199
transform 1 0 2876 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_2109
timestamp 1711653199
transform 1 0 2868 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1711653199
transform 1 0 3300 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2111
timestamp 1711653199
transform 1 0 3204 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1711653199
transform 1 0 3204 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1711653199
transform 1 0 3132 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1711653199
transform 1 0 3092 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2115
timestamp 1711653199
transform 1 0 3092 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1711653199
transform 1 0 3068 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1711653199
transform 1 0 3068 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1711653199
transform 1 0 3020 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1711653199
transform 1 0 3020 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1711653199
transform 1 0 2948 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1711653199
transform 1 0 2948 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1711653199
transform 1 0 2924 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1711653199
transform 1 0 2916 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1711653199
transform 1 0 2732 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1711653199
transform 1 0 2732 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1711653199
transform 1 0 2476 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1711653199
transform 1 0 2476 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1711653199
transform 1 0 2428 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1711653199
transform 1 0 2284 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1711653199
transform 1 0 2252 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1711653199
transform 1 0 2188 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1711653199
transform 1 0 2188 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1711653199
transform 1 0 2172 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1711653199
transform 1 0 2052 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1711653199
transform 1 0 2036 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1711653199
transform 1 0 2028 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1711653199
transform 1 0 1804 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2138
timestamp 1711653199
transform 1 0 1764 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1711653199
transform 1 0 1676 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1711653199
transform 1 0 1580 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1711653199
transform 1 0 1564 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1711653199
transform 1 0 1564 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1711653199
transform 1 0 1420 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1711653199
transform 1 0 1420 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1711653199
transform 1 0 1348 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1711653199
transform 1 0 1172 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1711653199
transform 1 0 1172 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1711653199
transform 1 0 1124 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1711653199
transform 1 0 964 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1711653199
transform 1 0 964 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1711653199
transform 1 0 916 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1711653199
transform 1 0 564 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_2153
timestamp 1711653199
transform 1 0 564 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1711653199
transform 1 0 540 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1711653199
transform 1 0 516 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1711653199
transform 1 0 516 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1711653199
transform 1 0 484 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1711653199
transform 1 0 484 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2159
timestamp 1711653199
transform 1 0 452 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2160
timestamp 1711653199
transform 1 0 452 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1711653199
transform 1 0 444 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2162
timestamp 1711653199
transform 1 0 444 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2163
timestamp 1711653199
transform 1 0 436 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1711653199
transform 1 0 436 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1711653199
transform 1 0 164 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1711653199
transform 1 0 164 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_2167
timestamp 1711653199
transform 1 0 124 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2168
timestamp 1711653199
transform 1 0 116 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2169
timestamp 1711653199
transform 1 0 108 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_2170
timestamp 1711653199
transform 1 0 2988 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2171
timestamp 1711653199
transform 1 0 2892 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1711653199
transform 1 0 2884 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1711653199
transform 1 0 2884 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2174
timestamp 1711653199
transform 1 0 2884 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2175
timestamp 1711653199
transform 1 0 2852 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2176
timestamp 1711653199
transform 1 0 2276 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1711653199
transform 1 0 2276 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2178
timestamp 1711653199
transform 1 0 2244 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2179
timestamp 1711653199
transform 1 0 1916 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2180
timestamp 1711653199
transform 1 0 1916 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_2181
timestamp 1711653199
transform 1 0 1844 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1711653199
transform 1 0 1772 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1711653199
transform 1 0 1724 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1711653199
transform 1 0 1636 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1711653199
transform 1 0 1636 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_2186
timestamp 1711653199
transform 1 0 1572 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1711653199
transform 1 0 1556 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1711653199
transform 1 0 1396 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2189
timestamp 1711653199
transform 1 0 1204 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1711653199
transform 1 0 1084 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1711653199
transform 1 0 948 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2192
timestamp 1711653199
transform 1 0 948 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2193
timestamp 1711653199
transform 1 0 828 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2194
timestamp 1711653199
transform 1 0 3356 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2195
timestamp 1711653199
transform 1 0 3260 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_2196
timestamp 1711653199
transform 1 0 3260 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1711653199
transform 1 0 3132 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2198
timestamp 1711653199
transform 1 0 3116 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2199
timestamp 1711653199
transform 1 0 3100 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_2200
timestamp 1711653199
transform 1 0 2868 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2201
timestamp 1711653199
transform 1 0 2860 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_2202
timestamp 1711653199
transform 1 0 2196 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2203
timestamp 1711653199
transform 1 0 1820 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2204
timestamp 1711653199
transform 1 0 1820 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_2205
timestamp 1711653199
transform 1 0 1748 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2206
timestamp 1711653199
transform 1 0 1740 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1711653199
transform 1 0 1700 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1711653199
transform 1 0 1700 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2209
timestamp 1711653199
transform 1 0 1500 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2210
timestamp 1711653199
transform 1 0 1500 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2211
timestamp 1711653199
transform 1 0 1356 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1711653199
transform 1 0 1180 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2213
timestamp 1711653199
transform 1 0 1100 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1711653199
transform 1 0 788 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1711653199
transform 1 0 404 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1711653199
transform 1 0 404 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_2217
timestamp 1711653199
transform 1 0 332 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2218
timestamp 1711653199
transform 1 0 236 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1711653199
transform 1 0 236 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1711653199
transform 1 0 180 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2221
timestamp 1711653199
transform 1 0 180 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1711653199
transform 1 0 3092 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2223
timestamp 1711653199
transform 1 0 2980 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1711653199
transform 1 0 2204 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1711653199
transform 1 0 2036 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1711653199
transform 1 0 1988 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2227
timestamp 1711653199
transform 1 0 1876 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1711653199
transform 1 0 1660 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2229
timestamp 1711653199
transform 1 0 1452 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2230
timestamp 1711653199
transform 1 0 1260 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2231
timestamp 1711653199
transform 1 0 1228 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2232
timestamp 1711653199
transform 1 0 1100 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1711653199
transform 1 0 460 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2234
timestamp 1711653199
transform 1 0 460 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1711653199
transform 1 0 420 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2236
timestamp 1711653199
transform 1 0 340 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2237
timestamp 1711653199
transform 1 0 244 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1711653199
transform 1 0 188 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1711653199
transform 1 0 188 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2240
timestamp 1711653199
transform 1 0 100 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2241
timestamp 1711653199
transform 1 0 2588 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_2242
timestamp 1711653199
transform 1 0 2444 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2243
timestamp 1711653199
transform 1 0 2404 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1711653199
transform 1 0 2276 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1711653199
transform 1 0 2244 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1711653199
transform 1 0 1676 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1711653199
transform 1 0 1676 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1711653199
transform 1 0 1620 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2249
timestamp 1711653199
transform 1 0 1428 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1711653199
transform 1 0 1404 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1711653199
transform 1 0 1364 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2252
timestamp 1711653199
transform 1 0 1308 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1711653199
transform 1 0 1308 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1711653199
transform 1 0 1196 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1711653199
transform 1 0 1188 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2256
timestamp 1711653199
transform 1 0 956 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1711653199
transform 1 0 900 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1711653199
transform 1 0 900 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1711653199
transform 1 0 620 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1711653199
transform 1 0 564 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2261
timestamp 1711653199
transform 1 0 532 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2262
timestamp 1711653199
transform 1 0 3148 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2263
timestamp 1711653199
transform 1 0 3132 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1711653199
transform 1 0 3076 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2265
timestamp 1711653199
transform 1 0 3076 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2266
timestamp 1711653199
transform 1 0 2940 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1711653199
transform 1 0 2884 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1711653199
transform 1 0 2884 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1711653199
transform 1 0 2812 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1711653199
transform 1 0 2772 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1711653199
transform 1 0 2772 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1711653199
transform 1 0 2652 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1711653199
transform 1 0 2652 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1711653199
transform 1 0 2436 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1711653199
transform 1 0 2404 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1711653199
transform 1 0 2404 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1711653199
transform 1 0 2364 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1711653199
transform 1 0 2308 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2279
timestamp 1711653199
transform 1 0 2156 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2280
timestamp 1711653199
transform 1 0 2820 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1711653199
transform 1 0 2820 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1711653199
transform 1 0 2796 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1711653199
transform 1 0 2740 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1711653199
transform 1 0 2740 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1711653199
transform 1 0 2636 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1711653199
transform 1 0 2636 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2287
timestamp 1711653199
transform 1 0 2596 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2288
timestamp 1711653199
transform 1 0 2596 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1711653199
transform 1 0 2180 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1711653199
transform 1 0 2172 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2291
timestamp 1711653199
transform 1 0 2132 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1711653199
transform 1 0 2132 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1711653199
transform 1 0 2092 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1711653199
transform 1 0 1972 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1711653199
transform 1 0 1972 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1711653199
transform 1 0 1852 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1711653199
transform 1 0 1700 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1711653199
transform 1 0 1628 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1711653199
transform 1 0 1044 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1711653199
transform 1 0 1044 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1711653199
transform 1 0 1036 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1711653199
transform 1 0 1004 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1711653199
transform 1 0 1004 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1711653199
transform 1 0 996 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1711653199
transform 1 0 988 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1711653199
transform 1 0 980 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1711653199
transform 1 0 956 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1711653199
transform 1 0 844 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1711653199
transform 1 0 844 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2310
timestamp 1711653199
transform 1 0 844 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1711653199
transform 1 0 796 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1711653199
transform 1 0 740 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2313
timestamp 1711653199
transform 1 0 636 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2314
timestamp 1711653199
transform 1 0 2828 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1711653199
transform 1 0 2596 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2316
timestamp 1711653199
transform 1 0 2596 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1711653199
transform 1 0 2548 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_2318
timestamp 1711653199
transform 1 0 2468 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1711653199
transform 1 0 2460 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1711653199
transform 1 0 2412 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2321
timestamp 1711653199
transform 1 0 2412 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_2322
timestamp 1711653199
transform 1 0 2380 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1711653199
transform 1 0 2180 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1711653199
transform 1 0 2172 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2325
timestamp 1711653199
transform 1 0 1884 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1711653199
transform 1 0 1836 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1711653199
transform 1 0 1796 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1711653199
transform 1 0 1772 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1711653199
transform 1 0 1772 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_2330
timestamp 1711653199
transform 1 0 1196 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1711653199
transform 1 0 1180 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1711653199
transform 1 0 996 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1711653199
transform 1 0 844 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1711653199
transform 1 0 844 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1711653199
transform 1 0 780 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1711653199
transform 1 0 764 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1711653199
transform 1 0 676 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1711653199
transform 1 0 3140 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2339
timestamp 1711653199
transform 1 0 3108 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1711653199
transform 1 0 3100 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_2341
timestamp 1711653199
transform 1 0 3052 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1711653199
transform 1 0 2252 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1711653199
transform 1 0 1988 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1711653199
transform 1 0 1988 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1711653199
transform 1 0 1972 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1711653199
transform 1 0 1972 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1711653199
transform 1 0 1804 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1711653199
transform 1 0 1716 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1711653199
transform 1 0 1716 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1711653199
transform 1 0 1604 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1711653199
transform 1 0 1604 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1711653199
transform 1 0 1508 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1711653199
transform 1 0 1508 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1711653199
transform 1 0 1340 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2355
timestamp 1711653199
transform 1 0 1004 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1711653199
transform 1 0 1004 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1711653199
transform 1 0 804 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_2358
timestamp 1711653199
transform 1 0 804 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2359
timestamp 1711653199
transform 1 0 780 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2360
timestamp 1711653199
transform 1 0 676 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2361
timestamp 1711653199
transform 1 0 524 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1711653199
transform 1 0 436 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1711653199
transform 1 0 436 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1711653199
transform 1 0 436 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2365
timestamp 1711653199
transform 1 0 348 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_2366
timestamp 1711653199
transform 1 0 2204 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1711653199
transform 1 0 2148 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1711653199
transform 1 0 1908 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2369
timestamp 1711653199
transform 1 0 1892 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2370
timestamp 1711653199
transform 1 0 1780 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1711653199
transform 1 0 1084 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1711653199
transform 1 0 1028 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2373
timestamp 1711653199
transform 1 0 972 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2374
timestamp 1711653199
transform 1 0 748 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1711653199
transform 1 0 676 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1711653199
transform 1 0 644 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2377
timestamp 1711653199
transform 1 0 644 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1711653199
transform 1 0 620 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2379
timestamp 1711653199
transform 1 0 588 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1711653199
transform 1 0 564 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_2381
timestamp 1711653199
transform 1 0 564 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1711653199
transform 1 0 3284 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1711653199
transform 1 0 3060 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1711653199
transform 1 0 2772 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1711653199
transform 1 0 2772 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1711653199
transform 1 0 2772 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_2387
timestamp 1711653199
transform 1 0 2668 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2388
timestamp 1711653199
transform 1 0 2660 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1711653199
transform 1 0 2412 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2390
timestamp 1711653199
transform 1 0 1748 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2391
timestamp 1711653199
transform 1 0 1748 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_2392
timestamp 1711653199
transform 1 0 1604 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2393
timestamp 1711653199
transform 1 0 1540 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1711653199
transform 1 0 1540 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1711653199
transform 1 0 1484 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2396
timestamp 1711653199
transform 1 0 1484 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1711653199
transform 1 0 1308 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1711653199
transform 1 0 812 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2399
timestamp 1711653199
transform 1 0 812 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1711653199
transform 1 0 556 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2401
timestamp 1711653199
transform 1 0 556 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_2402
timestamp 1711653199
transform 1 0 284 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2403
timestamp 1711653199
transform 1 0 212 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2404
timestamp 1711653199
transform 1 0 180 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2405
timestamp 1711653199
transform 1 0 172 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2406
timestamp 1711653199
transform 1 0 100 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2407
timestamp 1711653199
transform 1 0 68 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2408
timestamp 1711653199
transform 1 0 2508 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2409
timestamp 1711653199
transform 1 0 2468 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2410
timestamp 1711653199
transform 1 0 2412 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_2411
timestamp 1711653199
transform 1 0 2412 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2412
timestamp 1711653199
transform 1 0 2332 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1711653199
transform 1 0 2324 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2414
timestamp 1711653199
transform 1 0 1764 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_2415
timestamp 1711653199
transform 1 0 1764 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1711653199
transform 1 0 1708 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2417
timestamp 1711653199
transform 1 0 1708 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_2418
timestamp 1711653199
transform 1 0 1708 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2419
timestamp 1711653199
transform 1 0 1596 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2420
timestamp 1711653199
transform 1 0 1596 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1711653199
transform 1 0 1524 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2422
timestamp 1711653199
transform 1 0 1524 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1711653199
transform 1 0 1356 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1711653199
transform 1 0 1140 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2425
timestamp 1711653199
transform 1 0 1140 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2426
timestamp 1711653199
transform 1 0 1132 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2427
timestamp 1711653199
transform 1 0 1116 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2428
timestamp 1711653199
transform 1 0 780 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2429
timestamp 1711653199
transform 1 0 740 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2430
timestamp 1711653199
transform 1 0 604 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2431
timestamp 1711653199
transform 1 0 596 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1711653199
transform 1 0 588 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1711653199
transform 1 0 580 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1711653199
transform 1 0 324 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2435
timestamp 1711653199
transform 1 0 308 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2436
timestamp 1711653199
transform 1 0 292 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2437
timestamp 1711653199
transform 1 0 1268 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2438
timestamp 1711653199
transform 1 0 1108 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2439
timestamp 1711653199
transform 1 0 1052 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1711653199
transform 1 0 1004 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_2441
timestamp 1711653199
transform 1 0 1004 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2442
timestamp 1711653199
transform 1 0 956 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_2443
timestamp 1711653199
transform 1 0 956 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1711653199
transform 1 0 956 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2445
timestamp 1711653199
transform 1 0 852 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1711653199
transform 1 0 812 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2447
timestamp 1711653199
transform 1 0 668 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1711653199
transform 1 0 668 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2449
timestamp 1711653199
transform 1 0 660 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2450
timestamp 1711653199
transform 1 0 652 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2451
timestamp 1711653199
transform 1 0 452 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2452
timestamp 1711653199
transform 1 0 268 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2453
timestamp 1711653199
transform 1 0 260 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_2454
timestamp 1711653199
transform 1 0 3092 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2455
timestamp 1711653199
transform 1 0 3036 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1711653199
transform 1 0 3036 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1711653199
transform 1 0 2972 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2458
timestamp 1711653199
transform 1 0 3308 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2459
timestamp 1711653199
transform 1 0 3180 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2460
timestamp 1711653199
transform 1 0 3252 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_2461
timestamp 1711653199
transform 1 0 2956 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2462
timestamp 1711653199
transform 1 0 2396 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_2463
timestamp 1711653199
transform 1 0 3012 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2464
timestamp 1711653199
transform 1 0 2908 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2465
timestamp 1711653199
transform 1 0 2908 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_2466
timestamp 1711653199
transform 1 0 2732 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2467
timestamp 1711653199
transform 1 0 2196 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2468
timestamp 1711653199
transform 1 0 2172 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2469
timestamp 1711653199
transform 1 0 2036 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2470
timestamp 1711653199
transform 1 0 2036 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_2471
timestamp 1711653199
transform 1 0 1244 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_2472
timestamp 1711653199
transform 1 0 1212 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2473
timestamp 1711653199
transform 1 0 1148 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2474
timestamp 1711653199
transform 1 0 996 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2475
timestamp 1711653199
transform 1 0 2844 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2476
timestamp 1711653199
transform 1 0 2780 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2477
timestamp 1711653199
transform 1 0 2644 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2478
timestamp 1711653199
transform 1 0 2564 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1711653199
transform 1 0 2260 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1711653199
transform 1 0 2260 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1711653199
transform 1 0 2244 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2482
timestamp 1711653199
transform 1 0 1996 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2483
timestamp 1711653199
transform 1 0 1804 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1711653199
transform 1 0 3156 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1711653199
transform 1 0 3100 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1711653199
transform 1 0 3012 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2487
timestamp 1711653199
transform 1 0 2956 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1711653199
transform 1 0 2956 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1711653199
transform 1 0 2812 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_2490
timestamp 1711653199
transform 1 0 2812 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2491
timestamp 1711653199
transform 1 0 2748 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2492
timestamp 1711653199
transform 1 0 2724 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2493
timestamp 1711653199
transform 1 0 2724 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1711653199
transform 1 0 2268 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1711653199
transform 1 0 2900 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2496
timestamp 1711653199
transform 1 0 2788 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1711653199
transform 1 0 2788 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1711653199
transform 1 0 2084 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2499
timestamp 1711653199
transform 1 0 2076 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2500
timestamp 1711653199
transform 1 0 2012 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2501
timestamp 1711653199
transform 1 0 1996 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2502
timestamp 1711653199
transform 1 0 1332 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2503
timestamp 1711653199
transform 1 0 1332 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2504
timestamp 1711653199
transform 1 0 1332 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2505
timestamp 1711653199
transform 1 0 1292 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1711653199
transform 1 0 1244 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1711653199
transform 1 0 892 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1711653199
transform 1 0 892 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2509
timestamp 1711653199
transform 1 0 892 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1711653199
transform 1 0 828 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2511
timestamp 1711653199
transform 1 0 756 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1711653199
transform 1 0 716 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2513
timestamp 1711653199
transform 1 0 2612 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2514
timestamp 1711653199
transform 1 0 2308 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1711653199
transform 1 0 2836 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2516
timestamp 1711653199
transform 1 0 2748 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1711653199
transform 1 0 2700 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_2518
timestamp 1711653199
transform 1 0 3396 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1711653199
transform 1 0 3356 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1711653199
transform 1 0 3316 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1711653199
transform 1 0 2820 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1711653199
transform 1 0 2812 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1711653199
transform 1 0 2788 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1711653199
transform 1 0 2764 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_2525
timestamp 1711653199
transform 1 0 324 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1711653199
transform 1 0 284 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2527
timestamp 1711653199
transform 1 0 284 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1711653199
transform 1 0 284 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1711653199
transform 1 0 260 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1711653199
transform 1 0 260 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2531
timestamp 1711653199
transform 1 0 140 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_2532
timestamp 1711653199
transform 1 0 92 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1711653199
transform 1 0 2812 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1711653199
transform 1 0 2724 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2535
timestamp 1711653199
transform 1 0 2724 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2536
timestamp 1711653199
transform 1 0 2692 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1711653199
transform 1 0 2676 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_2538
timestamp 1711653199
transform 1 0 2636 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1711653199
transform 1 0 2636 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2540
timestamp 1711653199
transform 1 0 2628 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2541
timestamp 1711653199
transform 1 0 2628 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1711653199
transform 1 0 2604 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2543
timestamp 1711653199
transform 1 0 2188 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2544
timestamp 1711653199
transform 1 0 2156 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2545
timestamp 1711653199
transform 1 0 2028 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1711653199
transform 1 0 1748 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2547
timestamp 1711653199
transform 1 0 1132 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2548
timestamp 1711653199
transform 1 0 1132 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_2549
timestamp 1711653199
transform 1 0 924 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_2550
timestamp 1711653199
transform 1 0 3348 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1711653199
transform 1 0 3292 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_2552
timestamp 1711653199
transform 1 0 2964 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_2553
timestamp 1711653199
transform 1 0 2884 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_2554
timestamp 1711653199
transform 1 0 2820 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_2555
timestamp 1711653199
transform 1 0 2748 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_2556
timestamp 1711653199
transform 1 0 3116 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_2557
timestamp 1711653199
transform 1 0 3012 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1711653199
transform 1 0 2772 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_2559
timestamp 1711653199
transform 1 0 2708 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_2560
timestamp 1711653199
transform 1 0 3156 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2561
timestamp 1711653199
transform 1 0 3052 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2562
timestamp 1711653199
transform 1 0 3124 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2563
timestamp 1711653199
transform 1 0 3052 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2564
timestamp 1711653199
transform 1 0 2924 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2565
timestamp 1711653199
transform 1 0 2860 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_2566
timestamp 1711653199
transform 1 0 2764 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1711653199
transform 1 0 2692 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_2568
timestamp 1711653199
transform 1 0 2732 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1711653199
transform 1 0 2644 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2570
timestamp 1711653199
transform 1 0 3324 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2571
timestamp 1711653199
transform 1 0 3308 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2572
timestamp 1711653199
transform 1 0 3308 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2573
timestamp 1711653199
transform 1 0 3268 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2574
timestamp 1711653199
transform 1 0 3244 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2575
timestamp 1711653199
transform 1 0 3244 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2576
timestamp 1711653199
transform 1 0 3244 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2577
timestamp 1711653199
transform 1 0 3244 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2578
timestamp 1711653199
transform 1 0 3204 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_2579
timestamp 1711653199
transform 1 0 3204 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2580
timestamp 1711653199
transform 1 0 3140 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2581
timestamp 1711653199
transform 1 0 3140 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2582
timestamp 1711653199
transform 1 0 3068 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_2583
timestamp 1711653199
transform 1 0 3004 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2584
timestamp 1711653199
transform 1 0 2980 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_2585
timestamp 1711653199
transform 1 0 2980 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2586
timestamp 1711653199
transform 1 0 2932 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2587
timestamp 1711653199
transform 1 0 2932 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2588
timestamp 1711653199
transform 1 0 2812 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2589
timestamp 1711653199
transform 1 0 2812 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_2590
timestamp 1711653199
transform 1 0 2956 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_2591
timestamp 1711653199
transform 1 0 2892 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_2592
timestamp 1711653199
transform 1 0 2868 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2593
timestamp 1711653199
transform 1 0 2812 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_2594
timestamp 1711653199
transform 1 0 2908 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2595
timestamp 1711653199
transform 1 0 2828 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_2596
timestamp 1711653199
transform 1 0 3228 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2597
timestamp 1711653199
transform 1 0 3156 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_2598
timestamp 1711653199
transform 1 0 3108 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2599
timestamp 1711653199
transform 1 0 3028 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_2600
timestamp 1711653199
transform 1 0 2428 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_2601
timestamp 1711653199
transform 1 0 2284 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_2602
timestamp 1711653199
transform 1 0 2468 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_2603
timestamp 1711653199
transform 1 0 2388 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2604
timestamp 1711653199
transform 1 0 2356 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2605
timestamp 1711653199
transform 1 0 2236 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2606
timestamp 1711653199
transform 1 0 2676 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2607
timestamp 1711653199
transform 1 0 2604 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2608
timestamp 1711653199
transform 1 0 2300 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2609
timestamp 1711653199
transform 1 0 2076 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_2610
timestamp 1711653199
transform 1 0 1548 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2611
timestamp 1711653199
transform 1 0 1420 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_2612
timestamp 1711653199
transform 1 0 1660 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_2613
timestamp 1711653199
transform 1 0 1660 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_2614
timestamp 1711653199
transform 1 0 1612 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_2615
timestamp 1711653199
transform 1 0 1612 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_2616
timestamp 1711653199
transform 1 0 716 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2617
timestamp 1711653199
transform 1 0 604 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_2618
timestamp 1711653199
transform 1 0 980 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1711653199
transform 1 0 860 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1711653199
transform 1 0 220 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2621
timestamp 1711653199
transform 1 0 124 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_2622
timestamp 1711653199
transform 1 0 1132 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2623
timestamp 1711653199
transform 1 0 1092 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_2624
timestamp 1711653199
transform 1 0 1316 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2625
timestamp 1711653199
transform 1 0 1204 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2626
timestamp 1711653199
transform 1 0 1476 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2627
timestamp 1711653199
transform 1 0 1404 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_2628
timestamp 1711653199
transform 1 0 1676 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2629
timestamp 1711653199
transform 1 0 1564 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1711653199
transform 1 0 1924 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2631
timestamp 1711653199
transform 1 0 1836 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_2632
timestamp 1711653199
transform 1 0 3228 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2633
timestamp 1711653199
transform 1 0 3204 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2634
timestamp 1711653199
transform 1 0 3140 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2635
timestamp 1711653199
transform 1 0 3140 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2636
timestamp 1711653199
transform 1 0 2996 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2637
timestamp 1711653199
transform 1 0 2876 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_2638
timestamp 1711653199
transform 1 0 2876 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1711653199
transform 1 0 1828 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1711653199
transform 1 0 1828 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_2641
timestamp 1711653199
transform 1 0 1644 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1711653199
transform 1 0 1644 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2643
timestamp 1711653199
transform 1 0 1564 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2644
timestamp 1711653199
transform 1 0 1564 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2645
timestamp 1711653199
transform 1 0 1564 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_2646
timestamp 1711653199
transform 1 0 1556 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_2647
timestamp 1711653199
transform 1 0 1356 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1711653199
transform 1 0 780 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2649
timestamp 1711653199
transform 1 0 780 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_2650
timestamp 1711653199
transform 1 0 636 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2651
timestamp 1711653199
transform 1 0 468 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2652
timestamp 1711653199
transform 1 0 276 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2653
timestamp 1711653199
transform 1 0 220 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2654
timestamp 1711653199
transform 1 0 212 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2655
timestamp 1711653199
transform 1 0 3172 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2656
timestamp 1711653199
transform 1 0 3132 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_2657
timestamp 1711653199
transform 1 0 3132 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2658
timestamp 1711653199
transform 1 0 2964 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2659
timestamp 1711653199
transform 1 0 2732 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2660
timestamp 1711653199
transform 1 0 2308 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2661
timestamp 1711653199
transform 1 0 2308 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2662
timestamp 1711653199
transform 1 0 2284 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2663
timestamp 1711653199
transform 1 0 2124 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2664
timestamp 1711653199
transform 1 0 1668 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_2665
timestamp 1711653199
transform 1 0 1668 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2666
timestamp 1711653199
transform 1 0 1316 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2667
timestamp 1711653199
transform 1 0 748 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1711653199
transform 1 0 692 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1711653199
transform 1 0 588 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1711653199
transform 1 0 388 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2671
timestamp 1711653199
transform 1 0 236 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1711653199
transform 1 0 220 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2673
timestamp 1711653199
transform 1 0 196 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1711653199
transform 1 0 140 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1711653199
transform 1 0 140 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2676
timestamp 1711653199
transform 1 0 1644 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2677
timestamp 1711653199
transform 1 0 1548 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2678
timestamp 1711653199
transform 1 0 1748 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1711653199
transform 1 0 1628 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_2680
timestamp 1711653199
transform 1 0 3156 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2681
timestamp 1711653199
transform 1 0 3140 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_2682
timestamp 1711653199
transform 1 0 3100 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_2683
timestamp 1711653199
transform 1 0 3100 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2684
timestamp 1711653199
transform 1 0 2908 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2685
timestamp 1711653199
transform 1 0 2716 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1711653199
transform 1 0 3236 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1711653199
transform 1 0 3140 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2688
timestamp 1711653199
transform 1 0 3076 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_2689
timestamp 1711653199
transform 1 0 3076 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2690
timestamp 1711653199
transform 1 0 2452 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2691
timestamp 1711653199
transform 1 0 2444 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2692
timestamp 1711653199
transform 1 0 2380 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2693
timestamp 1711653199
transform 1 0 2364 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_2694
timestamp 1711653199
transform 1 0 3332 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2695
timestamp 1711653199
transform 1 0 3292 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1711653199
transform 1 0 3396 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2697
timestamp 1711653199
transform 1 0 3396 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1711653199
transform 1 0 3340 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_2699
timestamp 1711653199
transform 1 0 3340 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1711653199
transform 1 0 3244 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1711653199
transform 1 0 3164 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_2702
timestamp 1711653199
transform 1 0 3148 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2703
timestamp 1711653199
transform 1 0 3060 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1711653199
transform 1 0 3020 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2705
timestamp 1711653199
transform 1 0 2988 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1711653199
transform 1 0 2940 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2707
timestamp 1711653199
transform 1 0 2884 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1711653199
transform 1 0 2868 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2709
timestamp 1711653199
transform 1 0 2772 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1711653199
transform 1 0 2764 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2711
timestamp 1711653199
transform 1 0 2604 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1711653199
transform 1 0 2524 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2713
timestamp 1711653199
transform 1 0 2524 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_2714
timestamp 1711653199
transform 1 0 2444 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_2715
timestamp 1711653199
transform 1 0 2396 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1711653199
transform 1 0 1676 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2717
timestamp 1711653199
transform 1 0 1676 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2718
timestamp 1711653199
transform 1 0 1636 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_2719
timestamp 1711653199
transform 1 0 1636 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_2720
timestamp 1711653199
transform 1 0 1772 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2721
timestamp 1711653199
transform 1 0 1548 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2722
timestamp 1711653199
transform 1 0 2412 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2723
timestamp 1711653199
transform 1 0 1556 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_2724
timestamp 1711653199
transform 1 0 2780 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2725
timestamp 1711653199
transform 1 0 2732 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2726
timestamp 1711653199
transform 1 0 2724 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2727
timestamp 1711653199
transform 1 0 2580 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2728
timestamp 1711653199
transform 1 0 2476 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_2729
timestamp 1711653199
transform 1 0 2388 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2730
timestamp 1711653199
transform 1 0 1612 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2731
timestamp 1711653199
transform 1 0 1612 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2732
timestamp 1711653199
transform 1 0 1188 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2733
timestamp 1711653199
transform 1 0 2812 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2734
timestamp 1711653199
transform 1 0 2396 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2735
timestamp 1711653199
transform 1 0 2492 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2736
timestamp 1711653199
transform 1 0 2356 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_2737
timestamp 1711653199
transform 1 0 2340 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2738
timestamp 1711653199
transform 1 0 2284 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_2739
timestamp 1711653199
transform 1 0 2228 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1711653199
transform 1 0 2164 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2741
timestamp 1711653199
transform 1 0 2420 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2742
timestamp 1711653199
transform 1 0 2300 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2743
timestamp 1711653199
transform 1 0 3052 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2744
timestamp 1711653199
transform 1 0 2996 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2745
timestamp 1711653199
transform 1 0 2956 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2746
timestamp 1711653199
transform 1 0 2500 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2747
timestamp 1711653199
transform 1 0 2444 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_2748
timestamp 1711653199
transform 1 0 2500 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2749
timestamp 1711653199
transform 1 0 2300 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_2750
timestamp 1711653199
transform 1 0 2244 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2751
timestamp 1711653199
transform 1 0 2204 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_2752
timestamp 1711653199
transform 1 0 2172 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1711653199
transform 1 0 1884 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2754
timestamp 1711653199
transform 1 0 2348 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2755
timestamp 1711653199
transform 1 0 2140 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_2756
timestamp 1711653199
transform 1 0 2300 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2757
timestamp 1711653199
transform 1 0 2076 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_2758
timestamp 1711653199
transform 1 0 2036 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2759
timestamp 1711653199
transform 1 0 1972 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_2760
timestamp 1711653199
transform 1 0 2084 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2761
timestamp 1711653199
transform 1 0 1956 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2762
timestamp 1711653199
transform 1 0 2436 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2763
timestamp 1711653199
transform 1 0 2332 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_2764
timestamp 1711653199
transform 1 0 2532 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1711653199
transform 1 0 2420 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2766
timestamp 1711653199
transform 1 0 2468 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2767
timestamp 1711653199
transform 1 0 2420 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_2768
timestamp 1711653199
transform 1 0 2532 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2769
timestamp 1711653199
transform 1 0 2452 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2770
timestamp 1711653199
transform 1 0 2420 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2771
timestamp 1711653199
transform 1 0 3100 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2772
timestamp 1711653199
transform 1 0 2796 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2773
timestamp 1711653199
transform 1 0 2828 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2774
timestamp 1711653199
transform 1 0 2812 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2775
timestamp 1711653199
transform 1 0 2796 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2776
timestamp 1711653199
transform 1 0 2732 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_2777
timestamp 1711653199
transform 1 0 2732 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2778
timestamp 1711653199
transform 1 0 2628 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_2779
timestamp 1711653199
transform 1 0 2620 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2780
timestamp 1711653199
transform 1 0 2596 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2781
timestamp 1711653199
transform 1 0 2580 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2782
timestamp 1711653199
transform 1 0 2564 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2783
timestamp 1711653199
transform 1 0 2564 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2784
timestamp 1711653199
transform 1 0 2524 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2785
timestamp 1711653199
transform 1 0 2332 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_2786
timestamp 1711653199
transform 1 0 3076 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1711653199
transform 1 0 3076 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2788
timestamp 1711653199
transform 1 0 3044 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2789
timestamp 1711653199
transform 1 0 2948 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_2790
timestamp 1711653199
transform 1 0 2404 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2791
timestamp 1711653199
transform 1 0 1572 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_2792
timestamp 1711653199
transform 1 0 3196 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2793
timestamp 1711653199
transform 1 0 3084 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_2794
timestamp 1711653199
transform 1 0 3300 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2795
timestamp 1711653199
transform 1 0 3156 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2796
timestamp 1711653199
transform 1 0 3292 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2797
timestamp 1711653199
transform 1 0 3252 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2798
timestamp 1711653199
transform 1 0 3316 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2799
timestamp 1711653199
transform 1 0 3268 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2800
timestamp 1711653199
transform 1 0 1132 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2801
timestamp 1711653199
transform 1 0 612 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2802
timestamp 1711653199
transform 1 0 1140 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2803
timestamp 1711653199
transform 1 0 1020 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2804
timestamp 1711653199
transform 1 0 3180 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2805
timestamp 1711653199
transform 1 0 3012 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2806
timestamp 1711653199
transform 1 0 2972 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_2807
timestamp 1711653199
transform 1 0 2780 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2808
timestamp 1711653199
transform 1 0 2780 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2809
timestamp 1711653199
transform 1 0 2660 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2810
timestamp 1711653199
transform 1 0 2660 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2811
timestamp 1711653199
transform 1 0 2100 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2812
timestamp 1711653199
transform 1 0 2084 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_2813
timestamp 1711653199
transform 1 0 1724 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2814
timestamp 1711653199
transform 1 0 1268 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2815
timestamp 1711653199
transform 1 0 1268 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2816
timestamp 1711653199
transform 1 0 1196 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2817
timestamp 1711653199
transform 1 0 1132 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2818
timestamp 1711653199
transform 1 0 1020 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2819
timestamp 1711653199
transform 1 0 980 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_2820
timestamp 1711653199
transform 1 0 1012 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2821
timestamp 1711653199
transform 1 0 972 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2822
timestamp 1711653199
transform 1 0 948 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2823
timestamp 1711653199
transform 1 0 876 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2824
timestamp 1711653199
transform 1 0 780 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2825
timestamp 1711653199
transform 1 0 1124 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2826
timestamp 1711653199
transform 1 0 300 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2827
timestamp 1711653199
transform 1 0 1244 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2828
timestamp 1711653199
transform 1 0 1220 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2829
timestamp 1711653199
transform 1 0 1268 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2830
timestamp 1711653199
transform 1 0 1220 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2831
timestamp 1711653199
transform 1 0 252 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2832
timestamp 1711653199
transform 1 0 212 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_2833
timestamp 1711653199
transform 1 0 420 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2834
timestamp 1711653199
transform 1 0 332 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2835
timestamp 1711653199
transform 1 0 324 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_2836
timestamp 1711653199
transform 1 0 308 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_2837
timestamp 1711653199
transform 1 0 308 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2838
timestamp 1711653199
transform 1 0 532 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2839
timestamp 1711653199
transform 1 0 308 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_2840
timestamp 1711653199
transform 1 0 644 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2841
timestamp 1711653199
transform 1 0 572 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_2842
timestamp 1711653199
transform 1 0 692 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2843
timestamp 1711653199
transform 1 0 596 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2844
timestamp 1711653199
transform 1 0 524 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_2845
timestamp 1711653199
transform 1 0 724 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2846
timestamp 1711653199
transform 1 0 668 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_2847
timestamp 1711653199
transform 1 0 812 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2848
timestamp 1711653199
transform 1 0 740 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2849
timestamp 1711653199
transform 1 0 628 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_2850
timestamp 1711653199
transform 1 0 308 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2851
timestamp 1711653199
transform 1 0 268 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_2852
timestamp 1711653199
transform 1 0 348 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2853
timestamp 1711653199
transform 1 0 324 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_2854
timestamp 1711653199
transform 1 0 380 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2855
timestamp 1711653199
transform 1 0 372 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2856
timestamp 1711653199
transform 1 0 332 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2857
timestamp 1711653199
transform 1 0 164 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_2858
timestamp 1711653199
transform 1 0 444 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2859
timestamp 1711653199
transform 1 0 388 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_2860
timestamp 1711653199
transform 1 0 276 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2861
timestamp 1711653199
transform 1 0 148 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_2862
timestamp 1711653199
transform 1 0 324 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2863
timestamp 1711653199
transform 1 0 252 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2864
timestamp 1711653199
transform 1 0 220 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_2865
timestamp 1711653199
transform 1 0 2460 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2866
timestamp 1711653199
transform 1 0 2388 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2867
timestamp 1711653199
transform 1 0 2508 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2868
timestamp 1711653199
transform 1 0 2412 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1711653199
transform 1 0 2652 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2870
timestamp 1711653199
transform 1 0 2556 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2871
timestamp 1711653199
transform 1 0 2652 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2872
timestamp 1711653199
transform 1 0 620 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_2873
timestamp 1711653199
transform 1 0 532 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2874
timestamp 1711653199
transform 1 0 356 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_2875
timestamp 1711653199
transform 1 0 732 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2876
timestamp 1711653199
transform 1 0 652 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2877
timestamp 1711653199
transform 1 0 628 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_2878
timestamp 1711653199
transform 1 0 668 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2879
timestamp 1711653199
transform 1 0 548 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2880
timestamp 1711653199
transform 1 0 532 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2881
timestamp 1711653199
transform 1 0 460 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_2882
timestamp 1711653199
transform 1 0 356 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2883
timestamp 1711653199
transform 1 0 300 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_2884
timestamp 1711653199
transform 1 0 404 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2885
timestamp 1711653199
transform 1 0 380 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2886
timestamp 1711653199
transform 1 0 380 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_2887
timestamp 1711653199
transform 1 0 324 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2888
timestamp 1711653199
transform 1 0 284 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2889
timestamp 1711653199
transform 1 0 524 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2890
timestamp 1711653199
transform 1 0 428 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2891
timestamp 1711653199
transform 1 0 380 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_2892
timestamp 1711653199
transform 1 0 380 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_2893
timestamp 1711653199
transform 1 0 284 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2894
timestamp 1711653199
transform 1 0 132 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2895
timestamp 1711653199
transform 1 0 324 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2896
timestamp 1711653199
transform 1 0 284 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_2897
timestamp 1711653199
transform 1 0 2860 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2898
timestamp 1711653199
transform 1 0 2660 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2899
timestamp 1711653199
transform 1 0 2612 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_2900
timestamp 1711653199
transform 1 0 2740 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2901
timestamp 1711653199
transform 1 0 2532 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_2902
timestamp 1711653199
transform 1 0 2500 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2903
timestamp 1711653199
transform 1 0 1068 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_2904
timestamp 1711653199
transform 1 0 972 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2905
timestamp 1711653199
transform 1 0 908 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2906
timestamp 1711653199
transform 1 0 1276 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2907
timestamp 1711653199
transform 1 0 1108 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2908
timestamp 1711653199
transform 1 0 1092 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_2909
timestamp 1711653199
transform 1 0 1060 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_2910
timestamp 1711653199
transform 1 0 868 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2911
timestamp 1711653199
transform 1 0 284 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2912
timestamp 1711653199
transform 1 0 1252 0 1 35
box -3 -3 3 3
use M3_M2  M3_M2_2913
timestamp 1711653199
transform 1 0 956 0 1 35
box -3 -3 3 3
use M3_M2  M3_M2_2914
timestamp 1711653199
transform 1 0 1348 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2915
timestamp 1711653199
transform 1 0 1204 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_2916
timestamp 1711653199
transform 1 0 212 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2917
timestamp 1711653199
transform 1 0 180 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_2918
timestamp 1711653199
transform 1 0 460 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2919
timestamp 1711653199
transform 1 0 364 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_2920
timestamp 1711653199
transform 1 0 2972 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2921
timestamp 1711653199
transform 1 0 2796 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_2922
timestamp 1711653199
transform 1 0 3308 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2923
timestamp 1711653199
transform 1 0 2972 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_2924
timestamp 1711653199
transform 1 0 3380 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2925
timestamp 1711653199
transform 1 0 3340 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_2926
timestamp 1711653199
transform 1 0 3116 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2927
timestamp 1711653199
transform 1 0 3004 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_2928
timestamp 1711653199
transform 1 0 2460 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2929
timestamp 1711653199
transform 1 0 2332 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_2930
timestamp 1711653199
transform 1 0 2236 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1711653199
transform 1 0 2076 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_2932
timestamp 1711653199
transform 1 0 2660 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2933
timestamp 1711653199
transform 1 0 2572 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_2934
timestamp 1711653199
transform 1 0 2532 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_2935
timestamp 1711653199
transform 1 0 2460 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2936
timestamp 1711653199
transform 1 0 2396 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2937
timestamp 1711653199
transform 1 0 2324 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2938
timestamp 1711653199
transform 1 0 2260 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_2939
timestamp 1711653199
transform 1 0 2260 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2940
timestamp 1711653199
transform 1 0 2260 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_2941
timestamp 1711653199
transform 1 0 1900 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2942
timestamp 1711653199
transform 1 0 1484 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_2943
timestamp 1711653199
transform 1 0 2100 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2944
timestamp 1711653199
transform 1 0 2036 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2945
timestamp 1711653199
transform 1 0 1964 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_2946
timestamp 1711653199
transform 1 0 2084 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2947
timestamp 1711653199
transform 1 0 1852 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2948
timestamp 1711653199
transform 1 0 1852 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2949
timestamp 1711653199
transform 1 0 1748 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_2950
timestamp 1711653199
transform 1 0 2228 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_2951
timestamp 1711653199
transform 1 0 1924 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1711653199
transform 1 0 1892 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1711653199
transform 1 0 2340 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2954
timestamp 1711653199
transform 1 0 2324 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_2955
timestamp 1711653199
transform 1 0 2308 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2956
timestamp 1711653199
transform 1 0 2276 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_2957
timestamp 1711653199
transform 1 0 2428 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2958
timestamp 1711653199
transform 1 0 2300 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_2959
timestamp 1711653199
transform 1 0 2492 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2960
timestamp 1711653199
transform 1 0 2196 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_2961
timestamp 1711653199
transform 1 0 2324 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2962
timestamp 1711653199
transform 1 0 2132 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2963
timestamp 1711653199
transform 1 0 2508 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2964
timestamp 1711653199
transform 1 0 2356 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2965
timestamp 1711653199
transform 1 0 1764 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2966
timestamp 1711653199
transform 1 0 1684 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_2967
timestamp 1711653199
transform 1 0 1820 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2968
timestamp 1711653199
transform 1 0 1724 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_2969
timestamp 1711653199
transform 1 0 1916 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2970
timestamp 1711653199
transform 1 0 1844 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2971
timestamp 1711653199
transform 1 0 2556 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2972
timestamp 1711653199
transform 1 0 2396 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_2973
timestamp 1711653199
transform 1 0 2396 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2974
timestamp 1711653199
transform 1 0 1900 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2975
timestamp 1711653199
transform 1 0 2868 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2976
timestamp 1711653199
transform 1 0 2804 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2977
timestamp 1711653199
transform 1 0 2540 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_2978
timestamp 1711653199
transform 1 0 2644 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2979
timestamp 1711653199
transform 1 0 2548 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_2980
timestamp 1711653199
transform 1 0 2628 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2981
timestamp 1711653199
transform 1 0 2572 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2982
timestamp 1711653199
transform 1 0 2524 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_2983
timestamp 1711653199
transform 1 0 1868 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_2984
timestamp 1711653199
transform 1 0 1660 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2985
timestamp 1711653199
transform 1 0 1532 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_2986
timestamp 1711653199
transform 1 0 1956 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2987
timestamp 1711653199
transform 1 0 1892 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2988
timestamp 1711653199
transform 1 0 1636 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_2989
timestamp 1711653199
transform 1 0 2036 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2990
timestamp 1711653199
transform 1 0 1740 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2991
timestamp 1711653199
transform 1 0 1740 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2992
timestamp 1711653199
transform 1 0 788 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_2993
timestamp 1711653199
transform 1 0 1796 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2994
timestamp 1711653199
transform 1 0 1748 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_2995
timestamp 1711653199
transform 1 0 1724 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_2996
timestamp 1711653199
transform 1 0 1188 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_2997
timestamp 1711653199
transform 1 0 2788 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2998
timestamp 1711653199
transform 1 0 1772 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_2999
timestamp 1711653199
transform 1 0 3084 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3000
timestamp 1711653199
transform 1 0 2780 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3001
timestamp 1711653199
transform 1 0 2956 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3002
timestamp 1711653199
transform 1 0 2876 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3003
timestamp 1711653199
transform 1 0 2876 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3004
timestamp 1711653199
transform 1 0 2844 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3005
timestamp 1711653199
transform 1 0 2700 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3006
timestamp 1711653199
transform 1 0 2508 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3007
timestamp 1711653199
transform 1 0 2468 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3008
timestamp 1711653199
transform 1 0 2444 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3009
timestamp 1711653199
transform 1 0 3212 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3010
timestamp 1711653199
transform 1 0 3084 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3011
timestamp 1711653199
transform 1 0 3036 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3012
timestamp 1711653199
transform 1 0 3332 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3013
timestamp 1711653199
transform 1 0 3316 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3014
timestamp 1711653199
transform 1 0 3228 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3015
timestamp 1711653199
transform 1 0 3396 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3016
timestamp 1711653199
transform 1 0 3364 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3017
timestamp 1711653199
transform 1 0 3292 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3018
timestamp 1711653199
transform 1 0 3284 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3019
timestamp 1711653199
transform 1 0 3236 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3020
timestamp 1711653199
transform 1 0 1124 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_3021
timestamp 1711653199
transform 1 0 308 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_3022
timestamp 1711653199
transform 1 0 1244 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3023
timestamp 1711653199
transform 1 0 1148 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3024
timestamp 1711653199
transform 1 0 1180 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3025
timestamp 1711653199
transform 1 0 1092 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3026
timestamp 1711653199
transform 1 0 1060 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3027
timestamp 1711653199
transform 1 0 996 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3028
timestamp 1711653199
transform 1 0 940 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3029
timestamp 1711653199
transform 1 0 900 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3030
timestamp 1711653199
transform 1 0 876 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3031
timestamp 1711653199
transform 1 0 1124 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3032
timestamp 1711653199
transform 1 0 1004 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3033
timestamp 1711653199
transform 1 0 860 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3034
timestamp 1711653199
transform 1 0 892 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3035
timestamp 1711653199
transform 1 0 780 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3036
timestamp 1711653199
transform 1 0 1412 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3037
timestamp 1711653199
transform 1 0 1380 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3038
timestamp 1711653199
transform 1 0 1220 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3039
timestamp 1711653199
transform 1 0 1260 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3040
timestamp 1711653199
transform 1 0 1188 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3041
timestamp 1711653199
transform 1 0 308 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3042
timestamp 1711653199
transform 1 0 284 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3043
timestamp 1711653199
transform 1 0 428 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3044
timestamp 1711653199
transform 1 0 332 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3045
timestamp 1711653199
transform 1 0 748 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3046
timestamp 1711653199
transform 1 0 372 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3047
timestamp 1711653199
transform 1 0 780 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3048
timestamp 1711653199
transform 1 0 748 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3049
timestamp 1711653199
transform 1 0 796 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_3050
timestamp 1711653199
transform 1 0 780 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_3051
timestamp 1711653199
transform 1 0 732 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3052
timestamp 1711653199
transform 1 0 628 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3053
timestamp 1711653199
transform 1 0 980 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3054
timestamp 1711653199
transform 1 0 788 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3055
timestamp 1711653199
transform 1 0 772 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3056
timestamp 1711653199
transform 1 0 692 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3057
timestamp 1711653199
transform 1 0 684 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3058
timestamp 1711653199
transform 1 0 612 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3059
timestamp 1711653199
transform 1 0 380 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3060
timestamp 1711653199
transform 1 0 204 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_3061
timestamp 1711653199
transform 1 0 444 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3062
timestamp 1711653199
transform 1 0 420 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3063
timestamp 1711653199
transform 1 0 468 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3064
timestamp 1711653199
transform 1 0 420 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1711653199
transform 1 0 348 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3066
timestamp 1711653199
transform 1 0 580 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3067
timestamp 1711653199
transform 1 0 484 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3068
timestamp 1711653199
transform 1 0 2036 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3069
timestamp 1711653199
transform 1 0 2004 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1711653199
transform 1 0 2012 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3071
timestamp 1711653199
transform 1 0 1852 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3072
timestamp 1711653199
transform 1 0 2108 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3073
timestamp 1711653199
transform 1 0 2004 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3074
timestamp 1711653199
transform 1 0 2004 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3075
timestamp 1711653199
transform 1 0 1820 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3076
timestamp 1711653199
transform 1 0 1860 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3077
timestamp 1711653199
transform 1 0 1724 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1711653199
transform 1 0 1628 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3079
timestamp 1711653199
transform 1 0 2188 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3080
timestamp 1711653199
transform 1 0 2036 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3081
timestamp 1711653199
transform 1 0 2060 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3082
timestamp 1711653199
transform 1 0 2012 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3083
timestamp 1711653199
transform 1 0 2116 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3084
timestamp 1711653199
transform 1 0 1956 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3085
timestamp 1711653199
transform 1 0 1908 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3086
timestamp 1711653199
transform 1 0 2028 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3087
timestamp 1711653199
transform 1 0 1700 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3088
timestamp 1711653199
transform 1 0 1700 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_3089
timestamp 1711653199
transform 1 0 1668 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3090
timestamp 1711653199
transform 1 0 2332 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3091
timestamp 1711653199
transform 1 0 2228 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3092
timestamp 1711653199
transform 1 0 2172 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3093
timestamp 1711653199
transform 1 0 2284 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1711653199
transform 1 0 2204 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3095
timestamp 1711653199
transform 1 0 1484 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3096
timestamp 1711653199
transform 1 0 1452 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3097
timestamp 1711653199
transform 1 0 1724 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3098
timestamp 1711653199
transform 1 0 1412 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3099
timestamp 1711653199
transform 1 0 1452 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3100
timestamp 1711653199
transform 1 0 1412 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3101
timestamp 1711653199
transform 1 0 1428 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3102
timestamp 1711653199
transform 1 0 1124 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3103
timestamp 1711653199
transform 1 0 1116 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3104
timestamp 1711653199
transform 1 0 996 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3105
timestamp 1711653199
transform 1 0 2308 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1711653199
transform 1 0 2228 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3107
timestamp 1711653199
transform 1 0 1532 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3108
timestamp 1711653199
transform 1 0 1532 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3109
timestamp 1711653199
transform 1 0 1020 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3110
timestamp 1711653199
transform 1 0 1020 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3111
timestamp 1711653199
transform 1 0 948 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_3112
timestamp 1711653199
transform 1 0 900 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_3113
timestamp 1711653199
transform 1 0 900 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1711653199
transform 1 0 1364 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3115
timestamp 1711653199
transform 1 0 1308 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3116
timestamp 1711653199
transform 1 0 972 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_3117
timestamp 1711653199
transform 1 0 972 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3118
timestamp 1711653199
transform 1 0 956 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_3119
timestamp 1711653199
transform 1 0 1028 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3120
timestamp 1711653199
transform 1 0 1004 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3121
timestamp 1711653199
transform 1 0 948 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3122
timestamp 1711653199
transform 1 0 940 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3123
timestamp 1711653199
transform 1 0 708 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3124
timestamp 1711653199
transform 1 0 700 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3125
timestamp 1711653199
transform 1 0 684 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1711653199
transform 1 0 684 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3127
timestamp 1711653199
transform 1 0 668 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3128
timestamp 1711653199
transform 1 0 628 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3129
timestamp 1711653199
transform 1 0 1348 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3130
timestamp 1711653199
transform 1 0 1220 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_3131
timestamp 1711653199
transform 1 0 3204 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3132
timestamp 1711653199
transform 1 0 3196 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3133
timestamp 1711653199
transform 1 0 3076 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3134
timestamp 1711653199
transform 1 0 2956 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_3135
timestamp 1711653199
transform 1 0 2756 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3136
timestamp 1711653199
transform 1 0 2716 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3137
timestamp 1711653199
transform 1 0 1300 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3138
timestamp 1711653199
transform 1 0 1300 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_3139
timestamp 1711653199
transform 1 0 1236 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3140
timestamp 1711653199
transform 1 0 1228 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_3141
timestamp 1711653199
transform 1 0 1188 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_3142
timestamp 1711653199
transform 1 0 1436 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3143
timestamp 1711653199
transform 1 0 1324 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3144
timestamp 1711653199
transform 1 0 1268 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3145
timestamp 1711653199
transform 1 0 1244 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3146
timestamp 1711653199
transform 1 0 1212 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3147
timestamp 1711653199
transform 1 0 1196 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3148
timestamp 1711653199
transform 1 0 1492 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3149
timestamp 1711653199
transform 1 0 1388 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3150
timestamp 1711653199
transform 1 0 1276 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3151
timestamp 1711653199
transform 1 0 1244 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3152
timestamp 1711653199
transform 1 0 1180 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_3153
timestamp 1711653199
transform 1 0 860 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3154
timestamp 1711653199
transform 1 0 820 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3155
timestamp 1711653199
transform 1 0 804 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_3156
timestamp 1711653199
transform 1 0 1244 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3157
timestamp 1711653199
transform 1 0 836 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3158
timestamp 1711653199
transform 1 0 836 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3159
timestamp 1711653199
transform 1 0 628 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3160
timestamp 1711653199
transform 1 0 548 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3161
timestamp 1711653199
transform 1 0 548 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3162
timestamp 1711653199
transform 1 0 524 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3163
timestamp 1711653199
transform 1 0 492 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3164
timestamp 1711653199
transform 1 0 492 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3165
timestamp 1711653199
transform 1 0 1820 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3166
timestamp 1711653199
transform 1 0 1724 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3167
timestamp 1711653199
transform 1 0 2028 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3168
timestamp 1711653199
transform 1 0 1796 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3169
timestamp 1711653199
transform 1 0 2044 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3170
timestamp 1711653199
transform 1 0 1964 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3171
timestamp 1711653199
transform 1 0 1972 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3172
timestamp 1711653199
transform 1 0 1932 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3173
timestamp 1711653199
transform 1 0 1844 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3174
timestamp 1711653199
transform 1 0 1932 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3175
timestamp 1711653199
transform 1 0 1916 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3176
timestamp 1711653199
transform 1 0 1884 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3177
timestamp 1711653199
transform 1 0 1868 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3178
timestamp 1711653199
transform 1 0 1164 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3179
timestamp 1711653199
transform 1 0 1140 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3180
timestamp 1711653199
transform 1 0 2228 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3181
timestamp 1711653199
transform 1 0 2036 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3182
timestamp 1711653199
transform 1 0 1996 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3183
timestamp 1711653199
transform 1 0 1996 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3184
timestamp 1711653199
transform 1 0 1628 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3185
timestamp 1711653199
transform 1 0 812 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3186
timestamp 1711653199
transform 1 0 1988 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3187
timestamp 1711653199
transform 1 0 1876 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3188
timestamp 1711653199
transform 1 0 1876 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3189
timestamp 1711653199
transform 1 0 1836 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3190
timestamp 1711653199
transform 1 0 1836 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3191
timestamp 1711653199
transform 1 0 1700 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3192
timestamp 1711653199
transform 1 0 1700 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3193
timestamp 1711653199
transform 1 0 1644 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_3194
timestamp 1711653199
transform 1 0 1868 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3195
timestamp 1711653199
transform 1 0 1436 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3196
timestamp 1711653199
transform 1 0 1436 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3197
timestamp 1711653199
transform 1 0 1020 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3198
timestamp 1711653199
transform 1 0 1020 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3199
timestamp 1711653199
transform 1 0 876 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3200
timestamp 1711653199
transform 1 0 684 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3201
timestamp 1711653199
transform 1 0 564 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3202
timestamp 1711653199
transform 1 0 524 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3203
timestamp 1711653199
transform 1 0 524 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3204
timestamp 1711653199
transform 1 0 2972 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3205
timestamp 1711653199
transform 1 0 2964 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3206
timestamp 1711653199
transform 1 0 2956 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3207
timestamp 1711653199
transform 1 0 2932 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3208
timestamp 1711653199
transform 1 0 2932 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_3209
timestamp 1711653199
transform 1 0 2908 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3210
timestamp 1711653199
transform 1 0 2844 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3211
timestamp 1711653199
transform 1 0 2844 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3212
timestamp 1711653199
transform 1 0 1988 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3213
timestamp 1711653199
transform 1 0 1988 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_3214
timestamp 1711653199
transform 1 0 1884 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3215
timestamp 1711653199
transform 1 0 2556 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3216
timestamp 1711653199
transform 1 0 2516 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3217
timestamp 1711653199
transform 1 0 2364 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3218
timestamp 1711653199
transform 1 0 2356 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3219
timestamp 1711653199
transform 1 0 2300 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3220
timestamp 1711653199
transform 1 0 2284 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3221
timestamp 1711653199
transform 1 0 2276 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3222
timestamp 1711653199
transform 1 0 2276 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3223
timestamp 1711653199
transform 1 0 2268 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3224
timestamp 1711653199
transform 1 0 2228 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3225
timestamp 1711653199
transform 1 0 2220 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3226
timestamp 1711653199
transform 1 0 2084 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_3227
timestamp 1711653199
transform 1 0 1932 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3228
timestamp 1711653199
transform 1 0 1764 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3229
timestamp 1711653199
transform 1 0 1692 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3230
timestamp 1711653199
transform 1 0 1444 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_3231
timestamp 1711653199
transform 1 0 1428 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3232
timestamp 1711653199
transform 1 0 1388 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3233
timestamp 1711653199
transform 1 0 1084 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_3234
timestamp 1711653199
transform 1 0 1524 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3235
timestamp 1711653199
transform 1 0 1412 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3236
timestamp 1711653199
transform 1 0 1444 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3237
timestamp 1711653199
transform 1 0 1428 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3238
timestamp 1711653199
transform 1 0 1668 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3239
timestamp 1711653199
transform 1 0 1572 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3240
timestamp 1711653199
transform 1 0 1572 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3241
timestamp 1711653199
transform 1 0 1388 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3242
timestamp 1711653199
transform 1 0 1404 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3243
timestamp 1711653199
transform 1 0 1284 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3244
timestamp 1711653199
transform 1 0 1284 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3245
timestamp 1711653199
transform 1 0 292 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_3246
timestamp 1711653199
transform 1 0 252 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3247
timestamp 1711653199
transform 1 0 212 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3248
timestamp 1711653199
transform 1 0 172 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3249
timestamp 1711653199
transform 1 0 308 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3250
timestamp 1711653199
transform 1 0 284 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3251
timestamp 1711653199
transform 1 0 476 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1711653199
transform 1 0 468 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3253
timestamp 1711653199
transform 1 0 412 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3254
timestamp 1711653199
transform 1 0 364 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_3255
timestamp 1711653199
transform 1 0 364 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3256
timestamp 1711653199
transform 1 0 356 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_3257
timestamp 1711653199
transform 1 0 300 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3258
timestamp 1711653199
transform 1 0 1340 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3259
timestamp 1711653199
transform 1 0 1316 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3260
timestamp 1711653199
transform 1 0 324 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3261
timestamp 1711653199
transform 1 0 124 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3262
timestamp 1711653199
transform 1 0 124 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3263
timestamp 1711653199
transform 1 0 76 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3264
timestamp 1711653199
transform 1 0 76 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_3265
timestamp 1711653199
transform 1 0 76 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3266
timestamp 1711653199
transform 1 0 636 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3267
timestamp 1711653199
transform 1 0 332 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3268
timestamp 1711653199
transform 1 0 316 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3269
timestamp 1711653199
transform 1 0 308 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3270
timestamp 1711653199
transform 1 0 300 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3271
timestamp 1711653199
transform 1 0 268 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3272
timestamp 1711653199
transform 1 0 268 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3273
timestamp 1711653199
transform 1 0 236 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_3274
timestamp 1711653199
transform 1 0 2244 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_3275
timestamp 1711653199
transform 1 0 1724 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_3276
timestamp 1711653199
transform 1 0 2868 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_3277
timestamp 1711653199
transform 1 0 2604 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_3278
timestamp 1711653199
transform 1 0 2580 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3279
timestamp 1711653199
transform 1 0 2324 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3280
timestamp 1711653199
transform 1 0 2324 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3281
timestamp 1711653199
transform 1 0 2324 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1711653199
transform 1 0 2180 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3283
timestamp 1711653199
transform 1 0 1428 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3284
timestamp 1711653199
transform 1 0 2212 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3285
timestamp 1711653199
transform 1 0 2148 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3286
timestamp 1711653199
transform 1 0 2140 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3287
timestamp 1711653199
transform 1 0 2124 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3288
timestamp 1711653199
transform 1 0 1940 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3289
timestamp 1711653199
transform 1 0 2252 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_3290
timestamp 1711653199
transform 1 0 2196 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_3291
timestamp 1711653199
transform 1 0 2172 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3292
timestamp 1711653199
transform 1 0 2108 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3293
timestamp 1711653199
transform 1 0 2044 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3294
timestamp 1711653199
transform 1 0 3060 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3295
timestamp 1711653199
transform 1 0 2972 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3296
timestamp 1711653199
transform 1 0 2972 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3297
timestamp 1711653199
transform 1 0 1652 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3298
timestamp 1711653199
transform 1 0 2748 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3299
timestamp 1711653199
transform 1 0 2708 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3300
timestamp 1711653199
transform 1 0 2684 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3301
timestamp 1711653199
transform 1 0 1684 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3302
timestamp 1711653199
transform 1 0 1668 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3303
timestamp 1711653199
transform 1 0 1628 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3304
timestamp 1711653199
transform 1 0 1684 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3305
timestamp 1711653199
transform 1 0 1500 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3306
timestamp 1711653199
transform 1 0 1500 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3307
timestamp 1711653199
transform 1 0 1484 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3308
timestamp 1711653199
transform 1 0 1436 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3309
timestamp 1711653199
transform 1 0 1412 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_3310
timestamp 1711653199
transform 1 0 3044 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3311
timestamp 1711653199
transform 1 0 3028 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3312
timestamp 1711653199
transform 1 0 2956 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3313
timestamp 1711653199
transform 1 0 2924 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3314
timestamp 1711653199
transform 1 0 2436 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3315
timestamp 1711653199
transform 1 0 2436 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3316
timestamp 1711653199
transform 1 0 2372 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3317
timestamp 1711653199
transform 1 0 3124 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3318
timestamp 1711653199
transform 1 0 3084 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3319
timestamp 1711653199
transform 1 0 3348 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3320
timestamp 1711653199
transform 1 0 3276 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3321
timestamp 1711653199
transform 1 0 3276 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3322
timestamp 1711653199
transform 1 0 3252 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3323
timestamp 1711653199
transform 1 0 3244 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3324
timestamp 1711653199
transform 1 0 3116 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3325
timestamp 1711653199
transform 1 0 2852 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3326
timestamp 1711653199
transform 1 0 3284 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3327
timestamp 1711653199
transform 1 0 3236 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3328
timestamp 1711653199
transform 1 0 3228 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3329
timestamp 1711653199
transform 1 0 3140 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_3330
timestamp 1711653199
transform 1 0 2988 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3331
timestamp 1711653199
transform 1 0 1524 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3332
timestamp 1711653199
transform 1 0 1492 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_3333
timestamp 1711653199
transform 1 0 1508 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3334
timestamp 1711653199
transform 1 0 1484 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3335
timestamp 1711653199
transform 1 0 1484 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3336
timestamp 1711653199
transform 1 0 1180 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3337
timestamp 1711653199
transform 1 0 2852 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3338
timestamp 1711653199
transform 1 0 2788 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3339
timestamp 1711653199
transform 1 0 2748 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3340
timestamp 1711653199
transform 1 0 2748 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3341
timestamp 1711653199
transform 1 0 1100 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3342
timestamp 1711653199
transform 1 0 1084 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3343
timestamp 1711653199
transform 1 0 1084 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3344
timestamp 1711653199
transform 1 0 1084 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3345
timestamp 1711653199
transform 1 0 1052 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3346
timestamp 1711653199
transform 1 0 1052 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3347
timestamp 1711653199
transform 1 0 916 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_3348
timestamp 1711653199
transform 1 0 1372 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_3349
timestamp 1711653199
transform 1 0 1164 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3350
timestamp 1711653199
transform 1 0 1164 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3351
timestamp 1711653199
transform 1 0 1164 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3352
timestamp 1711653199
transform 1 0 1124 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3353
timestamp 1711653199
transform 1 0 1076 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3354
timestamp 1711653199
transform 1 0 1436 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3355
timestamp 1711653199
transform 1 0 1332 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3356
timestamp 1711653199
transform 1 0 1332 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3357
timestamp 1711653199
transform 1 0 1180 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3358
timestamp 1711653199
transform 1 0 1140 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3359
timestamp 1711653199
transform 1 0 1140 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3360
timestamp 1711653199
transform 1 0 1100 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_3361
timestamp 1711653199
transform 1 0 1076 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3362
timestamp 1711653199
transform 1 0 1180 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3363
timestamp 1711653199
transform 1 0 1044 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3364
timestamp 1711653199
transform 1 0 964 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3365
timestamp 1711653199
transform 1 0 964 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3366
timestamp 1711653199
transform 1 0 916 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3367
timestamp 1711653199
transform 1 0 892 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3368
timestamp 1711653199
transform 1 0 892 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3369
timestamp 1711653199
transform 1 0 868 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3370
timestamp 1711653199
transform 1 0 852 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3371
timestamp 1711653199
transform 1 0 732 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3372
timestamp 1711653199
transform 1 0 588 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_3373
timestamp 1711653199
transform 1 0 1508 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3374
timestamp 1711653199
transform 1 0 540 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3375
timestamp 1711653199
transform 1 0 1340 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3376
timestamp 1711653199
transform 1 0 1068 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_3377
timestamp 1711653199
transform 1 0 1068 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3378
timestamp 1711653199
transform 1 0 932 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3379
timestamp 1711653199
transform 1 0 548 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3380
timestamp 1711653199
transform 1 0 540 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3381
timestamp 1711653199
transform 1 0 532 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3382
timestamp 1711653199
transform 1 0 524 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_3383
timestamp 1711653199
transform 1 0 500 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3384
timestamp 1711653199
transform 1 0 500 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3385
timestamp 1711653199
transform 1 0 468 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3386
timestamp 1711653199
transform 1 0 732 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_3387
timestamp 1711653199
transform 1 0 516 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3388
timestamp 1711653199
transform 1 0 516 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3389
timestamp 1711653199
transform 1 0 500 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3390
timestamp 1711653199
transform 1 0 388 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3391
timestamp 1711653199
transform 1 0 380 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3392
timestamp 1711653199
transform 1 0 1428 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3393
timestamp 1711653199
transform 1 0 1196 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3394
timestamp 1711653199
transform 1 0 1196 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3395
timestamp 1711653199
transform 1 0 876 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3396
timestamp 1711653199
transform 1 0 780 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3397
timestamp 1711653199
transform 1 0 772 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3398
timestamp 1711653199
transform 1 0 700 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3399
timestamp 1711653199
transform 1 0 700 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3400
timestamp 1711653199
transform 1 0 580 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3401
timestamp 1711653199
transform 1 0 564 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3402
timestamp 1711653199
transform 1 0 524 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3403
timestamp 1711653199
transform 1 0 572 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3404
timestamp 1711653199
transform 1 0 548 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3405
timestamp 1711653199
transform 1 0 484 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_3406
timestamp 1711653199
transform 1 0 484 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3407
timestamp 1711653199
transform 1 0 340 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3408
timestamp 1711653199
transform 1 0 340 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_3409
timestamp 1711653199
transform 1 0 252 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3410
timestamp 1711653199
transform 1 0 252 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3411
timestamp 1711653199
transform 1 0 236 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3412
timestamp 1711653199
transform 1 0 1572 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3413
timestamp 1711653199
transform 1 0 1540 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3414
timestamp 1711653199
transform 1 0 1668 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3415
timestamp 1711653199
transform 1 0 1588 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3416
timestamp 1711653199
transform 1 0 2396 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_3417
timestamp 1711653199
transform 1 0 2076 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_3418
timestamp 1711653199
transform 1 0 2076 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3419
timestamp 1711653199
transform 1 0 1732 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3420
timestamp 1711653199
transform 1 0 2460 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3421
timestamp 1711653199
transform 1 0 2380 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3422
timestamp 1711653199
transform 1 0 2668 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3423
timestamp 1711653199
transform 1 0 2388 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3424
timestamp 1711653199
transform 1 0 2684 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_3425
timestamp 1711653199
transform 1 0 788 0 1 75
box -3 -3 3 3
use M3_M2  M3_M2_3426
timestamp 1711653199
transform 1 0 716 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3427
timestamp 1711653199
transform 1 0 388 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3428
timestamp 1711653199
transform 1 0 700 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3429
timestamp 1711653199
transform 1 0 636 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3430
timestamp 1711653199
transform 1 0 676 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3431
timestamp 1711653199
transform 1 0 620 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3432
timestamp 1711653199
transform 1 0 324 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3433
timestamp 1711653199
transform 1 0 308 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3434
timestamp 1711653199
transform 1 0 484 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_3435
timestamp 1711653199
transform 1 0 332 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3436
timestamp 1711653199
transform 1 0 228 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_3437
timestamp 1711653199
transform 1 0 460 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3438
timestamp 1711653199
transform 1 0 404 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3439
timestamp 1711653199
transform 1 0 260 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3440
timestamp 1711653199
transform 1 0 188 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3441
timestamp 1711653199
transform 1 0 132 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3442
timestamp 1711653199
transform 1 0 332 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3443
timestamp 1711653199
transform 1 0 252 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3444
timestamp 1711653199
transform 1 0 180 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3445
timestamp 1711653199
transform 1 0 2572 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3446
timestamp 1711653199
transform 1 0 2484 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3447
timestamp 1711653199
transform 1 0 2820 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_3448
timestamp 1711653199
transform 1 0 2604 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_3449
timestamp 1711653199
transform 1 0 2556 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_3450
timestamp 1711653199
transform 1 0 1148 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_3451
timestamp 1711653199
transform 1 0 1108 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3452
timestamp 1711653199
transform 1 0 956 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3453
timestamp 1711653199
transform 1 0 916 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3454
timestamp 1711653199
transform 1 0 764 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3455
timestamp 1711653199
transform 1 0 996 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3456
timestamp 1711653199
transform 1 0 964 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3457
timestamp 1711653199
transform 1 0 932 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_3458
timestamp 1711653199
transform 1 0 940 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_3459
timestamp 1711653199
transform 1 0 364 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_3460
timestamp 1711653199
transform 1 0 1164 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_3461
timestamp 1711653199
transform 1 0 1020 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_3462
timestamp 1711653199
transform 1 0 1276 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3463
timestamp 1711653199
transform 1 0 1156 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_3464
timestamp 1711653199
transform 1 0 340 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3465
timestamp 1711653199
transform 1 0 276 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3466
timestamp 1711653199
transform 1 0 188 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3467
timestamp 1711653199
transform 1 0 3100 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3468
timestamp 1711653199
transform 1 0 2860 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3469
timestamp 1711653199
transform 1 0 3380 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3470
timestamp 1711653199
transform 1 0 3204 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3471
timestamp 1711653199
transform 1 0 2540 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3472
timestamp 1711653199
transform 1 0 2468 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3473
timestamp 1711653199
transform 1 0 2436 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3474
timestamp 1711653199
transform 1 0 2220 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3475
timestamp 1711653199
transform 1 0 2780 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3476
timestamp 1711653199
transform 1 0 2628 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3477
timestamp 1711653199
transform 1 0 2580 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3478
timestamp 1711653199
transform 1 0 2580 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_3479
timestamp 1711653199
transform 1 0 2580 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3480
timestamp 1711653199
transform 1 0 2564 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3481
timestamp 1711653199
transform 1 0 2564 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3482
timestamp 1711653199
transform 1 0 2532 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_3483
timestamp 1711653199
transform 1 0 2780 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3484
timestamp 1711653199
transform 1 0 2652 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3485
timestamp 1711653199
transform 1 0 2652 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3486
timestamp 1711653199
transform 1 0 2588 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3487
timestamp 1711653199
transform 1 0 2548 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3488
timestamp 1711653199
transform 1 0 2356 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3489
timestamp 1711653199
transform 1 0 2452 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3490
timestamp 1711653199
transform 1 0 2340 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3491
timestamp 1711653199
transform 1 0 2476 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_3492
timestamp 1711653199
transform 1 0 2164 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_3493
timestamp 1711653199
transform 1 0 2292 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3494
timestamp 1711653199
transform 1 0 2188 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3495
timestamp 1711653199
transform 1 0 2436 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3496
timestamp 1711653199
transform 1 0 2404 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3497
timestamp 1711653199
transform 1 0 2388 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3498
timestamp 1711653199
transform 1 0 2460 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3499
timestamp 1711653199
transform 1 0 2404 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_3500
timestamp 1711653199
transform 1 0 1788 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3501
timestamp 1711653199
transform 1 0 1428 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3502
timestamp 1711653199
transform 1 0 940 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3503
timestamp 1711653199
transform 1 0 1748 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3504
timestamp 1711653199
transform 1 0 1652 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3505
timestamp 1711653199
transform 1 0 1652 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3506
timestamp 1711653199
transform 1 0 1388 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3507
timestamp 1711653199
transform 1 0 1588 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3508
timestamp 1711653199
transform 1 0 1532 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3509
timestamp 1711653199
transform 1 0 1548 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3510
timestamp 1711653199
transform 1 0 1524 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3511
timestamp 1711653199
transform 1 0 1508 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3512
timestamp 1711653199
transform 1 0 1468 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3513
timestamp 1711653199
transform 1 0 1812 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_3514
timestamp 1711653199
transform 1 0 1532 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3515
timestamp 1711653199
transform 1 0 1388 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3516
timestamp 1711653199
transform 1 0 1404 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3517
timestamp 1711653199
transform 1 0 1108 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3518
timestamp 1711653199
transform 1 0 1508 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3519
timestamp 1711653199
transform 1 0 548 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3520
timestamp 1711653199
transform 1 0 500 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3521
timestamp 1711653199
transform 1 0 388 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_3522
timestamp 1711653199
transform 1 0 548 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3523
timestamp 1711653199
transform 1 0 244 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3524
timestamp 1711653199
transform 1 0 2068 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3525
timestamp 1711653199
transform 1 0 1964 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3526
timestamp 1711653199
transform 1 0 1956 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_3527
timestamp 1711653199
transform 1 0 1740 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3528
timestamp 1711653199
transform 1 0 1612 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3529
timestamp 1711653199
transform 1 0 1532 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_3530
timestamp 1711653199
transform 1 0 2236 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_3531
timestamp 1711653199
transform 1 0 1548 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_3532
timestamp 1711653199
transform 1 0 1500 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3533
timestamp 1711653199
transform 1 0 604 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_3534
timestamp 1711653199
transform 1 0 604 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_3535
timestamp 1711653199
transform 1 0 140 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3536
timestamp 1711653199
transform 1 0 1276 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3537
timestamp 1711653199
transform 1 0 212 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3538
timestamp 1711653199
transform 1 0 148 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_3539
timestamp 1711653199
transform 1 0 148 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_3540
timestamp 1711653199
transform 1 0 124 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3541
timestamp 1711653199
transform 1 0 100 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_3542
timestamp 1711653199
transform 1 0 172 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3543
timestamp 1711653199
transform 1 0 92 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_3544
timestamp 1711653199
transform 1 0 84 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3545
timestamp 1711653199
transform 1 0 76 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3546
timestamp 1711653199
transform 1 0 148 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3547
timestamp 1711653199
transform 1 0 92 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3548
timestamp 1711653199
transform 1 0 228 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3549
timestamp 1711653199
transform 1 0 172 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3550
timestamp 1711653199
transform 1 0 124 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_3551
timestamp 1711653199
transform 1 0 324 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3552
timestamp 1711653199
transform 1 0 164 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_3553
timestamp 1711653199
transform 1 0 2356 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3554
timestamp 1711653199
transform 1 0 2212 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3555
timestamp 1711653199
transform 1 0 2364 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3556
timestamp 1711653199
transform 1 0 2284 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3557
timestamp 1711653199
transform 1 0 2460 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3558
timestamp 1711653199
transform 1 0 2356 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3559
timestamp 1711653199
transform 1 0 2300 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3560
timestamp 1711653199
transform 1 0 2292 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_3561
timestamp 1711653199
transform 1 0 2412 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3562
timestamp 1711653199
transform 1 0 2380 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3563
timestamp 1711653199
transform 1 0 2380 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3564
timestamp 1711653199
transform 1 0 2324 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3565
timestamp 1711653199
transform 1 0 2324 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_3566
timestamp 1711653199
transform 1 0 2260 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3567
timestamp 1711653199
transform 1 0 3084 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3568
timestamp 1711653199
transform 1 0 2892 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3569
timestamp 1711653199
transform 1 0 2892 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_3570
timestamp 1711653199
transform 1 0 1612 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_3571
timestamp 1711653199
transform 1 0 1628 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3572
timestamp 1711653199
transform 1 0 1380 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3573
timestamp 1711653199
transform 1 0 1260 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3574
timestamp 1711653199
transform 1 0 3148 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3575
timestamp 1711653199
transform 1 0 3108 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3576
timestamp 1711653199
transform 1 0 3052 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3577
timestamp 1711653199
transform 1 0 3052 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3578
timestamp 1711653199
transform 1 0 3220 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3579
timestamp 1711653199
transform 1 0 3116 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3580
timestamp 1711653199
transform 1 0 3356 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3581
timestamp 1711653199
transform 1 0 3268 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3582
timestamp 1711653199
transform 1 0 3212 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3583
timestamp 1711653199
transform 1 0 3364 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3584
timestamp 1711653199
transform 1 0 3292 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3585
timestamp 1711653199
transform 1 0 3252 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_3586
timestamp 1711653199
transform 1 0 1372 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3587
timestamp 1711653199
transform 1 0 1340 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_3588
timestamp 1711653199
transform 1 0 1364 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3589
timestamp 1711653199
transform 1 0 1060 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3590
timestamp 1711653199
transform 1 0 964 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3591
timestamp 1711653199
transform 1 0 860 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3592
timestamp 1711653199
transform 1 0 1020 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3593
timestamp 1711653199
transform 1 0 932 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3594
timestamp 1711653199
transform 1 0 1932 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3595
timestamp 1711653199
transform 1 0 1580 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3596
timestamp 1711653199
transform 1 0 1580 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3597
timestamp 1711653199
transform 1 0 1348 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_3598
timestamp 1711653199
transform 1 0 1364 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3599
timestamp 1711653199
transform 1 0 1236 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3600
timestamp 1711653199
transform 1 0 1876 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3601
timestamp 1711653199
transform 1 0 1796 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_3602
timestamp 1711653199
transform 1 0 2060 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3603
timestamp 1711653199
transform 1 0 1836 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3604
timestamp 1711653199
transform 1 0 2652 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3605
timestamp 1711653199
transform 1 0 2636 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3606
timestamp 1711653199
transform 1 0 2012 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_3607
timestamp 1711653199
transform 1 0 2164 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3608
timestamp 1711653199
transform 1 0 2140 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3609
timestamp 1711653199
transform 1 0 1980 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3610
timestamp 1711653199
transform 1 0 1972 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3611
timestamp 1711653199
transform 1 0 1900 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_3612
timestamp 1711653199
transform 1 0 1876 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3613
timestamp 1711653199
transform 1 0 1876 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_3614
timestamp 1711653199
transform 1 0 1860 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_3615
timestamp 1711653199
transform 1 0 1860 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_3616
timestamp 1711653199
transform 1 0 2172 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3617
timestamp 1711653199
transform 1 0 1844 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_3618
timestamp 1711653199
transform 1 0 1820 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3619
timestamp 1711653199
transform 1 0 1772 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3620
timestamp 1711653199
transform 1 0 1772 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_3621
timestamp 1711653199
transform 1 0 1684 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_3622
timestamp 1711653199
transform 1 0 1812 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3623
timestamp 1711653199
transform 1 0 804 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_3624
timestamp 1711653199
transform 1 0 732 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3625
timestamp 1711653199
transform 1 0 700 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3626
timestamp 1711653199
transform 1 0 2244 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3627
timestamp 1711653199
transform 1 0 1940 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3628
timestamp 1711653199
transform 1 0 1492 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3629
timestamp 1711653199
transform 1 0 740 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3630
timestamp 1711653199
transform 1 0 1636 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_3631
timestamp 1711653199
transform 1 0 1548 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_3632
timestamp 1711653199
transform 1 0 1828 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3633
timestamp 1711653199
transform 1 0 1692 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3634
timestamp 1711653199
transform 1 0 1716 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_3635
timestamp 1711653199
transform 1 0 1492 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_3636
timestamp 1711653199
transform 1 0 1924 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3637
timestamp 1711653199
transform 1 0 1788 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3638
timestamp 1711653199
transform 1 0 2148 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_3639
timestamp 1711653199
transform 1 0 1980 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3640
timestamp 1711653199
transform 1 0 1980 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_3641
timestamp 1711653199
transform 1 0 1900 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3642
timestamp 1711653199
transform 1 0 1924 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_3643
timestamp 1711653199
transform 1 0 852 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_3644
timestamp 1711653199
transform 1 0 3188 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3645
timestamp 1711653199
transform 1 0 2908 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3646
timestamp 1711653199
transform 1 0 2884 0 1 35
box -3 -3 3 3
use M3_M2  M3_M2_3647
timestamp 1711653199
transform 1 0 2316 0 1 35
box -3 -3 3 3
use M3_M2  M3_M2_3648
timestamp 1711653199
transform 1 0 2308 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_3649
timestamp 1711653199
transform 1 0 900 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3650
timestamp 1711653199
transform 1 0 900 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_3651
timestamp 1711653199
transform 1 0 836 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_3652
timestamp 1711653199
transform 1 0 916 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3653
timestamp 1711653199
transform 1 0 844 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3654
timestamp 1711653199
transform 1 0 860 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3655
timestamp 1711653199
transform 1 0 732 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3656
timestamp 1711653199
transform 1 0 676 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3657
timestamp 1711653199
transform 1 0 1452 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3658
timestamp 1711653199
transform 1 0 852 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3659
timestamp 1711653199
transform 1 0 588 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3660
timestamp 1711653199
transform 1 0 2484 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3661
timestamp 1711653199
transform 1 0 2228 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3662
timestamp 1711653199
transform 1 0 2228 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3663
timestamp 1711653199
transform 1 0 2180 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3664
timestamp 1711653199
transform 1 0 2108 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_3665
timestamp 1711653199
transform 1 0 2108 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_3666
timestamp 1711653199
transform 1 0 1468 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_3667
timestamp 1711653199
transform 1 0 1468 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_3668
timestamp 1711653199
transform 1 0 1244 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3669
timestamp 1711653199
transform 1 0 1004 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3670
timestamp 1711653199
transform 1 0 1004 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3671
timestamp 1711653199
transform 1 0 988 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_3672
timestamp 1711653199
transform 1 0 964 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3673
timestamp 1711653199
transform 1 0 956 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3674
timestamp 1711653199
transform 1 0 956 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3675
timestamp 1711653199
transform 1 0 956 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3676
timestamp 1711653199
transform 1 0 940 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3677
timestamp 1711653199
transform 1 0 940 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3678
timestamp 1711653199
transform 1 0 916 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3679
timestamp 1711653199
transform 1 0 916 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3680
timestamp 1711653199
transform 1 0 900 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_3681
timestamp 1711653199
transform 1 0 900 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_3682
timestamp 1711653199
transform 1 0 1428 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3683
timestamp 1711653199
transform 1 0 660 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3684
timestamp 1711653199
transform 1 0 612 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3685
timestamp 1711653199
transform 1 0 580 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3686
timestamp 1711653199
transform 1 0 1700 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3687
timestamp 1711653199
transform 1 0 1668 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3688
timestamp 1711653199
transform 1 0 1492 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_3689
timestamp 1711653199
transform 1 0 1524 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3690
timestamp 1711653199
transform 1 0 1340 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3691
timestamp 1711653199
transform 1 0 2556 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3692
timestamp 1711653199
transform 1 0 1948 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_3693
timestamp 1711653199
transform 1 0 2892 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3694
timestamp 1711653199
transform 1 0 2836 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3695
timestamp 1711653199
transform 1 0 2532 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3696
timestamp 1711653199
transform 1 0 2068 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3697
timestamp 1711653199
transform 1 0 2004 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3698
timestamp 1711653199
transform 1 0 2004 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3699
timestamp 1711653199
transform 1 0 1884 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3700
timestamp 1711653199
transform 1 0 1828 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_3701
timestamp 1711653199
transform 1 0 1932 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3702
timestamp 1711653199
transform 1 0 1820 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3703
timestamp 1711653199
transform 1 0 2196 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_3704
timestamp 1711653199
transform 1 0 2060 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3705
timestamp 1711653199
transform 1 0 1812 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3706
timestamp 1711653199
transform 1 0 260 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3707
timestamp 1711653199
transform 1 0 252 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_3708
timestamp 1711653199
transform 1 0 204 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3709
timestamp 1711653199
transform 1 0 780 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_3710
timestamp 1711653199
transform 1 0 684 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_3711
timestamp 1711653199
transform 1 0 700 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3712
timestamp 1711653199
transform 1 0 596 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_3713
timestamp 1711653199
transform 1 0 524 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3714
timestamp 1711653199
transform 1 0 196 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_3715
timestamp 1711653199
transform 1 0 236 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3716
timestamp 1711653199
transform 1 0 196 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3717
timestamp 1711653199
transform 1 0 196 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3718
timestamp 1711653199
transform 1 0 164 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_3719
timestamp 1711653199
transform 1 0 1668 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3720
timestamp 1711653199
transform 1 0 524 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_3721
timestamp 1711653199
transform 1 0 2972 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3722
timestamp 1711653199
transform 1 0 1660 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3723
timestamp 1711653199
transform 1 0 1676 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3724
timestamp 1711653199
transform 1 0 1332 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3725
timestamp 1711653199
transform 1 0 3124 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_3726
timestamp 1711653199
transform 1 0 3020 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3727
timestamp 1711653199
transform 1 0 3236 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3728
timestamp 1711653199
transform 1 0 3116 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3729
timestamp 1711653199
transform 1 0 3220 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3730
timestamp 1711653199
transform 1 0 3156 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3731
timestamp 1711653199
transform 1 0 412 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3732
timestamp 1711653199
transform 1 0 300 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_3733
timestamp 1711653199
transform 1 0 852 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3734
timestamp 1711653199
transform 1 0 764 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3735
timestamp 1711653199
transform 1 0 1284 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3736
timestamp 1711653199
transform 1 0 844 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3737
timestamp 1711653199
transform 1 0 1500 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3738
timestamp 1711653199
transform 1 0 1492 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3739
timestamp 1711653199
transform 1 0 1468 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3740
timestamp 1711653199
transform 1 0 1452 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3741
timestamp 1711653199
transform 1 0 1284 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3742
timestamp 1711653199
transform 1 0 1284 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3743
timestamp 1711653199
transform 1 0 1252 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_3744
timestamp 1711653199
transform 1 0 540 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_3745
timestamp 1711653199
transform 1 0 524 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3746
timestamp 1711653199
transform 1 0 244 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3747
timestamp 1711653199
transform 1 0 236 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3748
timestamp 1711653199
transform 1 0 236 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3749
timestamp 1711653199
transform 1 0 236 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3750
timestamp 1711653199
transform 1 0 212 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3751
timestamp 1711653199
transform 1 0 204 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_3752
timestamp 1711653199
transform 1 0 156 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3753
timestamp 1711653199
transform 1 0 148 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_3754
timestamp 1711653199
transform 1 0 1580 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3755
timestamp 1711653199
transform 1 0 1276 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_3756
timestamp 1711653199
transform 1 0 1300 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3757
timestamp 1711653199
transform 1 0 1252 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3758
timestamp 1711653199
transform 1 0 796 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3759
timestamp 1711653199
transform 1 0 764 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3760
timestamp 1711653199
transform 1 0 900 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3761
timestamp 1711653199
transform 1 0 860 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_3762
timestamp 1711653199
transform 1 0 860 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3763
timestamp 1711653199
transform 1 0 380 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3764
timestamp 1711653199
transform 1 0 268 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3765
timestamp 1711653199
transform 1 0 1100 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3766
timestamp 1711653199
transform 1 0 948 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3767
timestamp 1711653199
transform 1 0 1932 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3768
timestamp 1711653199
transform 1 0 1524 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_3769
timestamp 1711653199
transform 1 0 1572 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3770
timestamp 1711653199
transform 1 0 1524 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3771
timestamp 1711653199
transform 1 0 1508 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_3772
timestamp 1711653199
transform 1 0 852 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3773
timestamp 1711653199
transform 1 0 820 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3774
timestamp 1711653199
transform 1 0 724 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3775
timestamp 1711653199
transform 1 0 676 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_3776
timestamp 1711653199
transform 1 0 2364 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3777
timestamp 1711653199
transform 1 0 2068 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_3778
timestamp 1711653199
transform 1 0 2068 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_3779
timestamp 1711653199
transform 1 0 1740 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3780
timestamp 1711653199
transform 1 0 1132 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3781
timestamp 1711653199
transform 1 0 1132 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_3782
timestamp 1711653199
transform 1 0 876 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3783
timestamp 1711653199
transform 1 0 812 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3784
timestamp 1711653199
transform 1 0 804 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_3785
timestamp 1711653199
transform 1 0 684 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3786
timestamp 1711653199
transform 1 0 684 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3787
timestamp 1711653199
transform 1 0 660 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3788
timestamp 1711653199
transform 1 0 660 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3789
timestamp 1711653199
transform 1 0 660 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3790
timestamp 1711653199
transform 1 0 532 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_3791
timestamp 1711653199
transform 1 0 516 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3792
timestamp 1711653199
transform 1 0 468 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3793
timestamp 1711653199
transform 1 0 444 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3794
timestamp 1711653199
transform 1 0 436 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_3795
timestamp 1711653199
transform 1 0 396 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3796
timestamp 1711653199
transform 1 0 388 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3797
timestamp 1711653199
transform 1 0 364 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_3798
timestamp 1711653199
transform 1 0 356 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_3799
timestamp 1711653199
transform 1 0 340 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_3800
timestamp 1711653199
transform 1 0 332 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3801
timestamp 1711653199
transform 1 0 300 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_3802
timestamp 1711653199
transform 1 0 300 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3803
timestamp 1711653199
transform 1 0 876 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3804
timestamp 1711653199
transform 1 0 860 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3805
timestamp 1711653199
transform 1 0 876 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3806
timestamp 1711653199
transform 1 0 852 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3807
timestamp 1711653199
transform 1 0 892 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3808
timestamp 1711653199
transform 1 0 844 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_3809
timestamp 1711653199
transform 1 0 1500 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3810
timestamp 1711653199
transform 1 0 1236 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_3811
timestamp 1711653199
transform 1 0 1572 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3812
timestamp 1711653199
transform 1 0 1412 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_3813
timestamp 1711653199
transform 1 0 1404 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3814
timestamp 1711653199
transform 1 0 692 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3815
timestamp 1711653199
transform 1 0 1684 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3816
timestamp 1711653199
transform 1 0 1572 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3817
timestamp 1711653199
transform 1 0 1468 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_3818
timestamp 1711653199
transform 1 0 2108 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3819
timestamp 1711653199
transform 1 0 1996 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_3820
timestamp 1711653199
transform 1 0 2076 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3821
timestamp 1711653199
transform 1 0 2028 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3822
timestamp 1711653199
transform 1 0 1940 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_3823
timestamp 1711653199
transform 1 0 2564 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3824
timestamp 1711653199
transform 1 0 2540 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_3825
timestamp 1711653199
transform 1 0 2588 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3826
timestamp 1711653199
transform 1 0 2460 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3827
timestamp 1711653199
transform 1 0 2476 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3828
timestamp 1711653199
transform 1 0 2468 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3829
timestamp 1711653199
transform 1 0 2380 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_3830
timestamp 1711653199
transform 1 0 2156 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3831
timestamp 1711653199
transform 1 0 2516 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3832
timestamp 1711653199
transform 1 0 2460 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3833
timestamp 1711653199
transform 1 0 2356 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_3834
timestamp 1711653199
transform 1 0 2356 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_3835
timestamp 1711653199
transform 1 0 2588 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3836
timestamp 1711653199
transform 1 0 2508 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3837
timestamp 1711653199
transform 1 0 2404 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3838
timestamp 1711653199
transform 1 0 2060 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3839
timestamp 1711653199
transform 1 0 1988 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3840
timestamp 1711653199
transform 1 0 2164 0 1 25
box -3 -3 3 3
use M3_M2  M3_M2_3841
timestamp 1711653199
transform 1 0 2036 0 1 25
box -3 -3 3 3
use M3_M2  M3_M2_3842
timestamp 1711653199
transform 1 0 2060 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_3843
timestamp 1711653199
transform 1 0 1804 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_3844
timestamp 1711653199
transform 1 0 1604 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3845
timestamp 1711653199
transform 1 0 1460 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_3846
timestamp 1711653199
transform 1 0 1476 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3847
timestamp 1711653199
transform 1 0 124 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_3848
timestamp 1711653199
transform 1 0 308 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3849
timestamp 1711653199
transform 1 0 164 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_3850
timestamp 1711653199
transform 1 0 164 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3851
timestamp 1711653199
transform 1 0 100 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3852
timestamp 1711653199
transform 1 0 2884 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3853
timestamp 1711653199
transform 1 0 1644 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_3854
timestamp 1711653199
transform 1 0 3068 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3855
timestamp 1711653199
transform 1 0 2908 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3856
timestamp 1711653199
transform 1 0 3084 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3857
timestamp 1711653199
transform 1 0 3044 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_3858
timestamp 1711653199
transform 1 0 3212 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3859
timestamp 1711653199
transform 1 0 3100 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_3860
timestamp 1711653199
transform 1 0 1380 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3861
timestamp 1711653199
transform 1 0 1228 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3862
timestamp 1711653199
transform 1 0 1228 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_3863
timestamp 1711653199
transform 1 0 1188 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_3864
timestamp 1711653199
transform 1 0 1404 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3865
timestamp 1711653199
transform 1 0 1004 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3866
timestamp 1711653199
transform 1 0 980 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_3867
timestamp 1711653199
transform 1 0 1740 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3868
timestamp 1711653199
transform 1 0 1532 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3869
timestamp 1711653199
transform 1 0 1324 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3870
timestamp 1711653199
transform 1 0 1116 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3871
timestamp 1711653199
transform 1 0 932 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_3872
timestamp 1711653199
transform 1 0 1372 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3873
timestamp 1711653199
transform 1 0 492 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_3874
timestamp 1711653199
transform 1 0 444 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3875
timestamp 1711653199
transform 1 0 372 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_3876
timestamp 1711653199
transform 1 0 500 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3877
timestamp 1711653199
transform 1 0 220 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_3878
timestamp 1711653199
transform 1 0 2372 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_3879
timestamp 1711653199
transform 1 0 2188 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3880
timestamp 1711653199
transform 1 0 2156 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3881
timestamp 1711653199
transform 1 0 2100 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3882
timestamp 1711653199
transform 1 0 2068 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3883
timestamp 1711653199
transform 1 0 2068 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_3884
timestamp 1711653199
transform 1 0 2156 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3885
timestamp 1711653199
transform 1 0 2012 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_3886
timestamp 1711653199
transform 1 0 2748 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3887
timestamp 1711653199
transform 1 0 2540 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3888
timestamp 1711653199
transform 1 0 2484 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3889
timestamp 1711653199
transform 1 0 2412 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3890
timestamp 1711653199
transform 1 0 2388 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_3891
timestamp 1711653199
transform 1 0 2108 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3892
timestamp 1711653199
transform 1 0 2108 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3893
timestamp 1711653199
transform 1 0 2036 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3894
timestamp 1711653199
transform 1 0 2004 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_3895
timestamp 1711653199
transform 1 0 2332 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3896
timestamp 1711653199
transform 1 0 2140 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3897
timestamp 1711653199
transform 1 0 2132 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3898
timestamp 1711653199
transform 1 0 2060 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3899
timestamp 1711653199
transform 1 0 2060 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3900
timestamp 1711653199
transform 1 0 2012 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_3901
timestamp 1711653199
transform 1 0 1972 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3902
timestamp 1711653199
transform 1 0 1748 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3903
timestamp 1711653199
transform 1 0 2140 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_3904
timestamp 1711653199
transform 1 0 2084 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_3905
timestamp 1711653199
transform 1 0 2164 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3906
timestamp 1711653199
transform 1 0 2108 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_3907
timestamp 1711653199
transform 1 0 2244 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3908
timestamp 1711653199
transform 1 0 2156 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3909
timestamp 1711653199
transform 1 0 2156 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3910
timestamp 1711653199
transform 1 0 2092 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_3911
timestamp 1711653199
transform 1 0 2484 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_3912
timestamp 1711653199
transform 1 0 2228 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_3913
timestamp 1711653199
transform 1 0 2364 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3914
timestamp 1711653199
transform 1 0 2324 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_3915
timestamp 1711653199
transform 1 0 2196 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3916
timestamp 1711653199
transform 1 0 2100 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_3917
timestamp 1711653199
transform 1 0 2092 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_3918
timestamp 1711653199
transform 1 0 2444 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3919
timestamp 1711653199
transform 1 0 2412 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3920
timestamp 1711653199
transform 1 0 2396 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3921
timestamp 1711653199
transform 1 0 2396 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3922
timestamp 1711653199
transform 1 0 2156 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3923
timestamp 1711653199
transform 1 0 1908 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_3924
timestamp 1711653199
transform 1 0 2052 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3925
timestamp 1711653199
transform 1 0 2020 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3926
timestamp 1711653199
transform 1 0 1636 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_3927
timestamp 1711653199
transform 1 0 2276 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3928
timestamp 1711653199
transform 1 0 2068 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_3929
timestamp 1711653199
transform 1 0 2500 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3930
timestamp 1711653199
transform 1 0 2260 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_3931
timestamp 1711653199
transform 1 0 2292 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3932
timestamp 1711653199
transform 1 0 2260 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_3933
timestamp 1711653199
transform 1 0 2388 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3934
timestamp 1711653199
transform 1 0 2356 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3935
timestamp 1711653199
transform 1 0 2228 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3936
timestamp 1711653199
transform 1 0 2116 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_3937
timestamp 1711653199
transform 1 0 2588 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3938
timestamp 1711653199
transform 1 0 2540 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_3939
timestamp 1711653199
transform 1 0 2596 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3940
timestamp 1711653199
transform 1 0 2516 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3941
timestamp 1711653199
transform 1 0 2516 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3942
timestamp 1711653199
transform 1 0 2500 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_3943
timestamp 1711653199
transform 1 0 2484 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3944
timestamp 1711653199
transform 1 0 2164 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_3945
timestamp 1711653199
transform 1 0 3156 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3946
timestamp 1711653199
transform 1 0 2836 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3947
timestamp 1711653199
transform 1 0 2828 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_3948
timestamp 1711653199
transform 1 0 2780 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_3949
timestamp 1711653199
transform 1 0 2908 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3950
timestamp 1711653199
transform 1 0 2868 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3951
timestamp 1711653199
transform 1 0 2836 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_3952
timestamp 1711653199
transform 1 0 2716 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3953
timestamp 1711653199
transform 1 0 2652 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_3954
timestamp 1711653199
transform 1 0 2060 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3955
timestamp 1711653199
transform 1 0 2004 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_3956
timestamp 1711653199
transform 1 0 1988 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3957
timestamp 1711653199
transform 1 0 1924 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_3958
timestamp 1711653199
transform 1 0 2252 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3959
timestamp 1711653199
transform 1 0 2124 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_3960
timestamp 1711653199
transform 1 0 2108 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3961
timestamp 1711653199
transform 1 0 2028 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_3962
timestamp 1711653199
transform 1 0 2012 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3963
timestamp 1711653199
transform 1 0 1980 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_3964
timestamp 1711653199
transform 1 0 2012 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3965
timestamp 1711653199
transform 1 0 1964 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_3966
timestamp 1711653199
transform 1 0 1964 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3967
timestamp 1711653199
transform 1 0 1940 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_3968
timestamp 1711653199
transform 1 0 1940 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3969
timestamp 1711653199
transform 1 0 1908 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_3970
timestamp 1711653199
transform 1 0 2108 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3971
timestamp 1711653199
transform 1 0 2076 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_3972
timestamp 1711653199
transform 1 0 2172 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3973
timestamp 1711653199
transform 1 0 2116 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_3974
timestamp 1711653199
transform 1 0 2356 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3975
timestamp 1711653199
transform 1 0 2220 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3976
timestamp 1711653199
transform 1 0 2212 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_3977
timestamp 1711653199
transform 1 0 2140 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_3978
timestamp 1711653199
transform 1 0 2420 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3979
timestamp 1711653199
transform 1 0 2380 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3980
timestamp 1711653199
transform 1 0 2340 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3981
timestamp 1711653199
transform 1 0 2148 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_3982
timestamp 1711653199
transform 1 0 2148 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3983
timestamp 1711653199
transform 1 0 2116 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3984
timestamp 1711653199
transform 1 0 2100 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_3985
timestamp 1711653199
transform 1 0 2460 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3986
timestamp 1711653199
transform 1 0 2460 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3987
timestamp 1711653199
transform 1 0 2412 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_3988
timestamp 1711653199
transform 1 0 2236 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_3989
timestamp 1711653199
transform 1 0 2228 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3990
timestamp 1711653199
transform 1 0 2092 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3991
timestamp 1711653199
transform 1 0 1964 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3992
timestamp 1711653199
transform 1 0 1964 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_3993
timestamp 1711653199
transform 1 0 1636 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3994
timestamp 1711653199
transform 1 0 1636 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_3995
timestamp 1711653199
transform 1 0 1636 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3996
timestamp 1711653199
transform 1 0 1612 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_3997
timestamp 1711653199
transform 1 0 1524 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_3998
timestamp 1711653199
transform 1 0 2276 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_3999
timestamp 1711653199
transform 1 0 2124 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4000
timestamp 1711653199
transform 1 0 2060 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4001
timestamp 1711653199
transform 1 0 1772 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4002
timestamp 1711653199
transform 1 0 1668 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4003
timestamp 1711653199
transform 1 0 1652 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4004
timestamp 1711653199
transform 1 0 1620 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4005
timestamp 1711653199
transform 1 0 2324 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4006
timestamp 1711653199
transform 1 0 2284 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4007
timestamp 1711653199
transform 1 0 2396 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4008
timestamp 1711653199
transform 1 0 2308 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4009
timestamp 1711653199
transform 1 0 2356 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4010
timestamp 1711653199
transform 1 0 2188 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4011
timestamp 1711653199
transform 1 0 2164 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4012
timestamp 1711653199
transform 1 0 2148 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4013
timestamp 1711653199
transform 1 0 2196 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4014
timestamp 1711653199
transform 1 0 2124 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4015
timestamp 1711653199
transform 1 0 2108 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4016
timestamp 1711653199
transform 1 0 2012 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4017
timestamp 1711653199
transform 1 0 1964 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4018
timestamp 1711653199
transform 1 0 1868 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4019
timestamp 1711653199
transform 1 0 1820 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4020
timestamp 1711653199
transform 1 0 1580 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4021
timestamp 1711653199
transform 1 0 1508 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4022
timestamp 1711653199
transform 1 0 1436 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4023
timestamp 1711653199
transform 1 0 1068 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4024
timestamp 1711653199
transform 1 0 1996 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4025
timestamp 1711653199
transform 1 0 1596 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4026
timestamp 1711653199
transform 1 0 1596 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4027
timestamp 1711653199
transform 1 0 1100 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4028
timestamp 1711653199
transform 1 0 1060 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4029
timestamp 1711653199
transform 1 0 756 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4030
timestamp 1711653199
transform 1 0 2100 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4031
timestamp 1711653199
transform 1 0 2044 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4032
timestamp 1711653199
transform 1 0 2044 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4033
timestamp 1711653199
transform 1 0 1956 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4034
timestamp 1711653199
transform 1 0 1956 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4035
timestamp 1711653199
transform 1 0 1900 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4036
timestamp 1711653199
transform 1 0 1788 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4037
timestamp 1711653199
transform 1 0 1684 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4038
timestamp 1711653199
transform 1 0 2020 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4039
timestamp 1711653199
transform 1 0 1796 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4040
timestamp 1711653199
transform 1 0 1796 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4041
timestamp 1711653199
transform 1 0 1772 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4042
timestamp 1711653199
transform 1 0 1900 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4043
timestamp 1711653199
transform 1 0 1780 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4044
timestamp 1711653199
transform 1 0 1908 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4045
timestamp 1711653199
transform 1 0 1868 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4046
timestamp 1711653199
transform 1 0 1964 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4047
timestamp 1711653199
transform 1 0 1924 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4048
timestamp 1711653199
transform 1 0 1900 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4049
timestamp 1711653199
transform 1 0 1892 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4050
timestamp 1711653199
transform 1 0 2068 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4051
timestamp 1711653199
transform 1 0 2068 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_4052
timestamp 1711653199
transform 1 0 2044 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4053
timestamp 1711653199
transform 1 0 2044 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4054
timestamp 1711653199
transform 1 0 2044 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_4055
timestamp 1711653199
transform 1 0 1908 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4056
timestamp 1711653199
transform 1 0 2348 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4057
timestamp 1711653199
transform 1 0 2156 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4058
timestamp 1711653199
transform 1 0 2068 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4059
timestamp 1711653199
transform 1 0 1996 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4060
timestamp 1711653199
transform 1 0 1812 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4061
timestamp 1711653199
transform 1 0 1500 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4062
timestamp 1711653199
transform 1 0 1500 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4063
timestamp 1711653199
transform 1 0 1340 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_4064
timestamp 1711653199
transform 1 0 1340 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4065
timestamp 1711653199
transform 1 0 1340 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_4066
timestamp 1711653199
transform 1 0 1308 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_4067
timestamp 1711653199
transform 1 0 1308 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_4068
timestamp 1711653199
transform 1 0 564 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4069
timestamp 1711653199
transform 1 0 420 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4070
timestamp 1711653199
transform 1 0 420 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4071
timestamp 1711653199
transform 1 0 404 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_4072
timestamp 1711653199
transform 1 0 396 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4073
timestamp 1711653199
transform 1 0 308 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_4074
timestamp 1711653199
transform 1 0 268 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_4075
timestamp 1711653199
transform 1 0 252 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_4076
timestamp 1711653199
transform 1 0 1892 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4077
timestamp 1711653199
transform 1 0 1804 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4078
timestamp 1711653199
transform 1 0 1804 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4079
timestamp 1711653199
transform 1 0 1788 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4080
timestamp 1711653199
transform 1 0 1740 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4081
timestamp 1711653199
transform 1 0 1724 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_4082
timestamp 1711653199
transform 1 0 932 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_4083
timestamp 1711653199
transform 1 0 908 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4084
timestamp 1711653199
transform 1 0 684 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4085
timestamp 1711653199
transform 1 0 2372 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4086
timestamp 1711653199
transform 1 0 2332 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4087
timestamp 1711653199
transform 1 0 2332 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4088
timestamp 1711653199
transform 1 0 2220 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4089
timestamp 1711653199
transform 1 0 1940 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4090
timestamp 1711653199
transform 1 0 1876 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4091
timestamp 1711653199
transform 1 0 1836 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4092
timestamp 1711653199
transform 1 0 884 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4093
timestamp 1711653199
transform 1 0 868 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4094
timestamp 1711653199
transform 1 0 860 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4095
timestamp 1711653199
transform 1 0 2164 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4096
timestamp 1711653199
transform 1 0 1996 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_4097
timestamp 1711653199
transform 1 0 2068 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4098
timestamp 1711653199
transform 1 0 2004 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4099
timestamp 1711653199
transform 1 0 2756 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4100
timestamp 1711653199
transform 1 0 2692 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_4101
timestamp 1711653199
transform 1 0 2676 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4102
timestamp 1711653199
transform 1 0 2676 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_4103
timestamp 1711653199
transform 1 0 2332 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4104
timestamp 1711653199
transform 1 0 2332 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_4105
timestamp 1711653199
transform 1 0 2180 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4106
timestamp 1711653199
transform 1 0 2156 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4107
timestamp 1711653199
transform 1 0 2076 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4108
timestamp 1711653199
transform 1 0 1948 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4109
timestamp 1711653199
transform 1 0 1796 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4110
timestamp 1711653199
transform 1 0 1740 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4111
timestamp 1711653199
transform 1 0 1196 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4112
timestamp 1711653199
transform 1 0 1004 0 1 675
box -3 -3 3 3
use M3_M2  M3_M2_4113
timestamp 1711653199
transform 1 0 1004 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4114
timestamp 1711653199
transform 1 0 716 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4115
timestamp 1711653199
transform 1 0 708 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_4116
timestamp 1711653199
transform 1 0 580 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4117
timestamp 1711653199
transform 1 0 564 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4118
timestamp 1711653199
transform 1 0 500 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4119
timestamp 1711653199
transform 1 0 3012 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4120
timestamp 1711653199
transform 1 0 3012 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4121
timestamp 1711653199
transform 1 0 3012 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_4122
timestamp 1711653199
transform 1 0 2868 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_4123
timestamp 1711653199
transform 1 0 2828 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_4124
timestamp 1711653199
transform 1 0 2140 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4125
timestamp 1711653199
transform 1 0 2140 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_4126
timestamp 1711653199
transform 1 0 2028 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_4127
timestamp 1711653199
transform 1 0 1308 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4128
timestamp 1711653199
transform 1 0 1300 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4129
timestamp 1711653199
transform 1 0 1260 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4130
timestamp 1711653199
transform 1 0 956 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4131
timestamp 1711653199
transform 1 0 884 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4132
timestamp 1711653199
transform 1 0 884 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4133
timestamp 1711653199
transform 1 0 844 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4134
timestamp 1711653199
transform 1 0 780 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_4135
timestamp 1711653199
transform 1 0 780 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4136
timestamp 1711653199
transform 1 0 724 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_4137
timestamp 1711653199
transform 1 0 2156 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4138
timestamp 1711653199
transform 1 0 2132 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4139
timestamp 1711653199
transform 1 0 2300 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4140
timestamp 1711653199
transform 1 0 1812 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4141
timestamp 1711653199
transform 1 0 1772 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4142
timestamp 1711653199
transform 1 0 1700 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4143
timestamp 1711653199
transform 1 0 1684 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4144
timestamp 1711653199
transform 1 0 900 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4145
timestamp 1711653199
transform 1 0 2836 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4146
timestamp 1711653199
transform 1 0 2596 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4147
timestamp 1711653199
transform 1 0 2396 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_4148
timestamp 1711653199
transform 1 0 2268 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4149
timestamp 1711653199
transform 1 0 2244 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4150
timestamp 1711653199
transform 1 0 1844 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4151
timestamp 1711653199
transform 1 0 1796 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4152
timestamp 1711653199
transform 1 0 1260 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4153
timestamp 1711653199
transform 1 0 1252 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4154
timestamp 1711653199
transform 1 0 1004 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4155
timestamp 1711653199
transform 1 0 1884 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4156
timestamp 1711653199
transform 1 0 1820 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4157
timestamp 1711653199
transform 1 0 1580 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4158
timestamp 1711653199
transform 1 0 1524 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4159
timestamp 1711653199
transform 1 0 1604 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4160
timestamp 1711653199
transform 1 0 1540 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4161
timestamp 1711653199
transform 1 0 1708 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4162
timestamp 1711653199
transform 1 0 1548 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4163
timestamp 1711653199
transform 1 0 1724 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4164
timestamp 1711653199
transform 1 0 1676 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4165
timestamp 1711653199
transform 1 0 1900 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4166
timestamp 1711653199
transform 1 0 1748 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4167
timestamp 1711653199
transform 1 0 2228 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4168
timestamp 1711653199
transform 1 0 1964 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4169
timestamp 1711653199
transform 1 0 1924 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4170
timestamp 1711653199
transform 1 0 1892 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4171
timestamp 1711653199
transform 1 0 1628 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4172
timestamp 1711653199
transform 1 0 1612 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4173
timestamp 1711653199
transform 1 0 1300 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_4174
timestamp 1711653199
transform 1 0 1300 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4175
timestamp 1711653199
transform 1 0 1012 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_4176
timestamp 1711653199
transform 1 0 1012 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4177
timestamp 1711653199
transform 1 0 596 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4178
timestamp 1711653199
transform 1 0 596 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_4179
timestamp 1711653199
transform 1 0 348 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4180
timestamp 1711653199
transform 1 0 348 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4181
timestamp 1711653199
transform 1 0 260 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4182
timestamp 1711653199
transform 1 0 260 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4183
timestamp 1711653199
transform 1 0 236 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4184
timestamp 1711653199
transform 1 0 228 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4185
timestamp 1711653199
transform 1 0 108 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4186
timestamp 1711653199
transform 1 0 92 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4187
timestamp 1711653199
transform 1 0 1900 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4188
timestamp 1711653199
transform 1 0 1716 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_4189
timestamp 1711653199
transform 1 0 1684 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4190
timestamp 1711653199
transform 1 0 1628 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_4191
timestamp 1711653199
transform 1 0 1716 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4192
timestamp 1711653199
transform 1 0 1684 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4193
timestamp 1711653199
transform 1 0 1596 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4194
timestamp 1711653199
transform 1 0 1588 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4195
timestamp 1711653199
transform 1 0 1588 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4196
timestamp 1711653199
transform 1 0 1516 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4197
timestamp 1711653199
transform 1 0 1372 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4198
timestamp 1711653199
transform 1 0 1708 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_4199
timestamp 1711653199
transform 1 0 1708 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4200
timestamp 1711653199
transform 1 0 1636 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4201
timestamp 1711653199
transform 1 0 1596 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_4202
timestamp 1711653199
transform 1 0 1660 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4203
timestamp 1711653199
transform 1 0 1548 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4204
timestamp 1711653199
transform 1 0 1156 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4205
timestamp 1711653199
transform 1 0 604 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_4206
timestamp 1711653199
transform 1 0 2484 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4207
timestamp 1711653199
transform 1 0 2452 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4208
timestamp 1711653199
transform 1 0 2356 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4209
timestamp 1711653199
transform 1 0 2348 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4210
timestamp 1711653199
transform 1 0 2132 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4211
timestamp 1711653199
transform 1 0 2132 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4212
timestamp 1711653199
transform 1 0 2100 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4213
timestamp 1711653199
transform 1 0 2092 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4214
timestamp 1711653199
transform 1 0 2044 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4215
timestamp 1711653199
transform 1 0 1620 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4216
timestamp 1711653199
transform 1 0 1612 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4217
timestamp 1711653199
transform 1 0 1588 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4218
timestamp 1711653199
transform 1 0 1436 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4219
timestamp 1711653199
transform 1 0 1436 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4220
timestamp 1711653199
transform 1 0 1108 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_4221
timestamp 1711653199
transform 1 0 1964 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4222
timestamp 1711653199
transform 1 0 1796 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_4223
timestamp 1711653199
transform 1 0 2028 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4224
timestamp 1711653199
transform 1 0 1988 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4225
timestamp 1711653199
transform 1 0 2444 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4226
timestamp 1711653199
transform 1 0 2420 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4227
timestamp 1711653199
transform 1 0 2420 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_4228
timestamp 1711653199
transform 1 0 1716 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4229
timestamp 1711653199
transform 1 0 1716 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4230
timestamp 1711653199
transform 1 0 1572 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4231
timestamp 1711653199
transform 1 0 1524 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4232
timestamp 1711653199
transform 1 0 1276 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_4233
timestamp 1711653199
transform 1 0 812 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4234
timestamp 1711653199
transform 1 0 2932 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4235
timestamp 1711653199
transform 1 0 2932 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4236
timestamp 1711653199
transform 1 0 2804 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4237
timestamp 1711653199
transform 1 0 2636 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4238
timestamp 1711653199
transform 1 0 2404 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4239
timestamp 1711653199
transform 1 0 1772 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4240
timestamp 1711653199
transform 1 0 1772 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4241
timestamp 1711653199
transform 1 0 1556 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4242
timestamp 1711653199
transform 1 0 1500 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4243
timestamp 1711653199
transform 1 0 1844 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4244
timestamp 1711653199
transform 1 0 1836 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4245
timestamp 1711653199
transform 1 0 1812 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4246
timestamp 1711653199
transform 1 0 1812 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4247
timestamp 1711653199
transform 1 0 1732 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4248
timestamp 1711653199
transform 1 0 1692 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4249
timestamp 1711653199
transform 1 0 1692 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4250
timestamp 1711653199
transform 1 0 1228 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4251
timestamp 1711653199
transform 1 0 1228 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4252
timestamp 1711653199
transform 1 0 812 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4253
timestamp 1711653199
transform 1 0 1300 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4254
timestamp 1711653199
transform 1 0 1260 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4255
timestamp 1711653199
transform 1 0 964 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4256
timestamp 1711653199
transform 1 0 772 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4257
timestamp 1711653199
transform 1 0 772 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4258
timestamp 1711653199
transform 1 0 668 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4259
timestamp 1711653199
transform 1 0 1572 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4260
timestamp 1711653199
transform 1 0 1324 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4261
timestamp 1711653199
transform 1 0 1612 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4262
timestamp 1711653199
transform 1 0 1548 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4263
timestamp 1711653199
transform 1 0 1836 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4264
timestamp 1711653199
transform 1 0 1836 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4265
timestamp 1711653199
transform 1 0 1708 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4266
timestamp 1711653199
transform 1 0 1300 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4267
timestamp 1711653199
transform 1 0 1300 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4268
timestamp 1711653199
transform 1 0 1284 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4269
timestamp 1711653199
transform 1 0 1268 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4270
timestamp 1711653199
transform 1 0 1156 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4271
timestamp 1711653199
transform 1 0 660 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4272
timestamp 1711653199
transform 1 0 660 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_4273
timestamp 1711653199
transform 1 0 404 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4274
timestamp 1711653199
transform 1 0 404 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4275
timestamp 1711653199
transform 1 0 340 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4276
timestamp 1711653199
transform 1 0 316 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_4277
timestamp 1711653199
transform 1 0 316 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4278
timestamp 1711653199
transform 1 0 316 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4279
timestamp 1711653199
transform 1 0 292 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4280
timestamp 1711653199
transform 1 0 292 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4281
timestamp 1711653199
transform 1 0 180 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4282
timestamp 1711653199
transform 1 0 164 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4283
timestamp 1711653199
transform 1 0 164 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4284
timestamp 1711653199
transform 1 0 1796 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4285
timestamp 1711653199
transform 1 0 1668 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4286
timestamp 1711653199
transform 1 0 1636 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4287
timestamp 1711653199
transform 1 0 1556 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4288
timestamp 1711653199
transform 1 0 1556 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_4289
timestamp 1711653199
transform 1 0 1548 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4290
timestamp 1711653199
transform 1 0 1644 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_4291
timestamp 1711653199
transform 1 0 1644 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4292
timestamp 1711653199
transform 1 0 1588 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4293
timestamp 1711653199
transform 1 0 1452 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_4294
timestamp 1711653199
transform 1 0 1340 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_4295
timestamp 1711653199
transform 1 0 1924 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4296
timestamp 1711653199
transform 1 0 1740 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4297
timestamp 1711653199
transform 1 0 1700 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4298
timestamp 1711653199
transform 1 0 1668 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_4299
timestamp 1711653199
transform 1 0 1660 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4300
timestamp 1711653199
transform 1 0 1628 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4301
timestamp 1711653199
transform 1 0 1516 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4302
timestamp 1711653199
transform 1 0 1244 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4303
timestamp 1711653199
transform 1 0 1052 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4304
timestamp 1711653199
transform 1 0 908 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4305
timestamp 1711653199
transform 1 0 1564 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4306
timestamp 1711653199
transform 1 0 1540 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4307
timestamp 1711653199
transform 1 0 1572 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4308
timestamp 1711653199
transform 1 0 1548 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_4309
timestamp 1711653199
transform 1 0 1820 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4310
timestamp 1711653199
transform 1 0 1668 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4311
timestamp 1711653199
transform 1 0 1924 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4312
timestamp 1711653199
transform 1 0 1828 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4313
timestamp 1711653199
transform 1 0 2348 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4314
timestamp 1711653199
transform 1 0 1500 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4315
timestamp 1711653199
transform 1 0 1500 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4316
timestamp 1711653199
transform 1 0 1484 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4317
timestamp 1711653199
transform 1 0 1228 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4318
timestamp 1711653199
transform 1 0 1220 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4319
timestamp 1711653199
transform 1 0 1116 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4320
timestamp 1711653199
transform 1 0 1116 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4321
timestamp 1711653199
transform 1 0 876 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4322
timestamp 1711653199
transform 1 0 2948 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4323
timestamp 1711653199
transform 1 0 2820 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4324
timestamp 1711653199
transform 1 0 2684 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4325
timestamp 1711653199
transform 1 0 2420 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4326
timestamp 1711653199
transform 1 0 1532 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4327
timestamp 1711653199
transform 1 0 1860 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4328
timestamp 1711653199
transform 1 0 1836 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_4329
timestamp 1711653199
transform 1 0 1796 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4330
timestamp 1711653199
transform 1 0 1620 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4331
timestamp 1711653199
transform 1 0 1620 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4332
timestamp 1711653199
transform 1 0 1604 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4333
timestamp 1711653199
transform 1 0 1604 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4334
timestamp 1711653199
transform 1 0 1604 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4335
timestamp 1711653199
transform 1 0 1548 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_4336
timestamp 1711653199
transform 1 0 1076 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4337
timestamp 1711653199
transform 1 0 1012 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4338
timestamp 1711653199
transform 1 0 1244 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4339
timestamp 1711653199
transform 1 0 972 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4340
timestamp 1711653199
transform 1 0 972 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4341
timestamp 1711653199
transform 1 0 660 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4342
timestamp 1711653199
transform 1 0 300 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4343
timestamp 1711653199
transform 1 0 2028 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4344
timestamp 1711653199
transform 1 0 1180 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4345
timestamp 1711653199
transform 1 0 1172 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4346
timestamp 1711653199
transform 1 0 1172 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4347
timestamp 1711653199
transform 1 0 1132 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4348
timestamp 1711653199
transform 1 0 1132 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4349
timestamp 1711653199
transform 1 0 2044 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4350
timestamp 1711653199
transform 1 0 1932 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4351
timestamp 1711653199
transform 1 0 2116 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4352
timestamp 1711653199
transform 1 0 2108 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4353
timestamp 1711653199
transform 1 0 2100 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4354
timestamp 1711653199
transform 1 0 2084 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_4355
timestamp 1711653199
transform 1 0 2084 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4356
timestamp 1711653199
transform 1 0 2060 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4357
timestamp 1711653199
transform 1 0 2060 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4358
timestamp 1711653199
transform 1 0 2044 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4359
timestamp 1711653199
transform 1 0 1948 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_4360
timestamp 1711653199
transform 1 0 1916 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4361
timestamp 1711653199
transform 1 0 1596 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4362
timestamp 1711653199
transform 1 0 1156 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4363
timestamp 1711653199
transform 1 0 2108 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4364
timestamp 1711653199
transform 1 0 2036 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4365
timestamp 1711653199
transform 1 0 1580 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4366
timestamp 1711653199
transform 1 0 1580 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4367
timestamp 1711653199
transform 1 0 756 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_4368
timestamp 1711653199
transform 1 0 2204 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4369
timestamp 1711653199
transform 1 0 2012 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_4370
timestamp 1711653199
transform 1 0 1860 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4371
timestamp 1711653199
transform 1 0 1644 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4372
timestamp 1711653199
transform 1 0 1644 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4373
timestamp 1711653199
transform 1 0 1044 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4374
timestamp 1711653199
transform 1 0 940 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4375
timestamp 1711653199
transform 1 0 1228 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4376
timestamp 1711653199
transform 1 0 1124 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4377
timestamp 1711653199
transform 1 0 876 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4378
timestamp 1711653199
transform 1 0 788 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4379
timestamp 1711653199
transform 1 0 740 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4380
timestamp 1711653199
transform 1 0 1908 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4381
timestamp 1711653199
transform 1 0 1876 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4382
timestamp 1711653199
transform 1 0 2036 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4383
timestamp 1711653199
transform 1 0 1956 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4384
timestamp 1711653199
transform 1 0 1908 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4385
timestamp 1711653199
transform 1 0 1908 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4386
timestamp 1711653199
transform 1 0 1732 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4387
timestamp 1711653199
transform 1 0 500 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4388
timestamp 1711653199
transform 1 0 372 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4389
timestamp 1711653199
transform 1 0 564 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4390
timestamp 1711653199
transform 1 0 452 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_4391
timestamp 1711653199
transform 1 0 604 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4392
timestamp 1711653199
transform 1 0 452 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_4393
timestamp 1711653199
transform 1 0 628 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4394
timestamp 1711653199
transform 1 0 604 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4395
timestamp 1711653199
transform 1 0 692 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4396
timestamp 1711653199
transform 1 0 668 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4397
timestamp 1711653199
transform 1 0 844 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4398
timestamp 1711653199
transform 1 0 676 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4399
timestamp 1711653199
transform 1 0 644 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4400
timestamp 1711653199
transform 1 0 628 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4401
timestamp 1711653199
transform 1 0 604 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4402
timestamp 1711653199
transform 1 0 668 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4403
timestamp 1711653199
transform 1 0 628 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_4404
timestamp 1711653199
transform 1 0 652 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_4405
timestamp 1711653199
transform 1 0 644 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4406
timestamp 1711653199
transform 1 0 1516 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4407
timestamp 1711653199
transform 1 0 732 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_4408
timestamp 1711653199
transform 1 0 732 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4409
timestamp 1711653199
transform 1 0 628 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4410
timestamp 1711653199
transform 1 0 588 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4411
timestamp 1711653199
transform 1 0 588 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_4412
timestamp 1711653199
transform 1 0 364 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4413
timestamp 1711653199
transform 1 0 620 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_4414
timestamp 1711653199
transform 1 0 556 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_4415
timestamp 1711653199
transform 1 0 2884 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_4416
timestamp 1711653199
transform 1 0 2820 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_4417
timestamp 1711653199
transform 1 0 2724 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_4418
timestamp 1711653199
transform 1 0 2580 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_4419
timestamp 1711653199
transform 1 0 2580 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_4420
timestamp 1711653199
transform 1 0 1964 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4421
timestamp 1711653199
transform 1 0 1852 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4422
timestamp 1711653199
transform 1 0 684 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4423
timestamp 1711653199
transform 1 0 628 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4424
timestamp 1711653199
transform 1 0 700 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4425
timestamp 1711653199
transform 1 0 636 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4426
timestamp 1711653199
transform 1 0 988 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4427
timestamp 1711653199
transform 1 0 708 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4428
timestamp 1711653199
transform 1 0 2324 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4429
timestamp 1711653199
transform 1 0 2252 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4430
timestamp 1711653199
transform 1 0 2244 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4431
timestamp 1711653199
transform 1 0 2212 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4432
timestamp 1711653199
transform 1 0 1996 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4433
timestamp 1711653199
transform 1 0 1996 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4434
timestamp 1711653199
transform 1 0 1900 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4435
timestamp 1711653199
transform 1 0 1596 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4436
timestamp 1711653199
transform 1 0 260 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4437
timestamp 1711653199
transform 1 0 124 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4438
timestamp 1711653199
transform 1 0 76 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4439
timestamp 1711653199
transform 1 0 76 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_4440
timestamp 1711653199
transform 1 0 188 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4441
timestamp 1711653199
transform 1 0 76 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_4442
timestamp 1711653199
transform 1 0 148 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4443
timestamp 1711653199
transform 1 0 108 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_4444
timestamp 1711653199
transform 1 0 228 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4445
timestamp 1711653199
transform 1 0 116 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4446
timestamp 1711653199
transform 1 0 228 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4447
timestamp 1711653199
transform 1 0 180 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4448
timestamp 1711653199
transform 1 0 348 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4449
timestamp 1711653199
transform 1 0 348 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4450
timestamp 1711653199
transform 1 0 316 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4451
timestamp 1711653199
transform 1 0 228 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4452
timestamp 1711653199
transform 1 0 172 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4453
timestamp 1711653199
transform 1 0 276 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4454
timestamp 1711653199
transform 1 0 244 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4455
timestamp 1711653199
transform 1 0 564 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4456
timestamp 1711653199
transform 1 0 548 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_4457
timestamp 1711653199
transform 1 0 428 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4458
timestamp 1711653199
transform 1 0 412 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4459
timestamp 1711653199
transform 1 0 236 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_4460
timestamp 1711653199
transform 1 0 228 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4461
timestamp 1711653199
transform 1 0 196 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4462
timestamp 1711653199
transform 1 0 196 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4463
timestamp 1711653199
transform 1 0 188 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4464
timestamp 1711653199
transform 1 0 172 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4465
timestamp 1711653199
transform 1 0 220 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_4466
timestamp 1711653199
transform 1 0 204 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4467
timestamp 1711653199
transform 1 0 188 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4468
timestamp 1711653199
transform 1 0 188 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_4469
timestamp 1711653199
transform 1 0 220 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4470
timestamp 1711653199
transform 1 0 188 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_4471
timestamp 1711653199
transform 1 0 252 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4472
timestamp 1711653199
transform 1 0 132 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4473
timestamp 1711653199
transform 1 0 212 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4474
timestamp 1711653199
transform 1 0 196 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_4475
timestamp 1711653199
transform 1 0 364 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4476
timestamp 1711653199
transform 1 0 340 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_4477
timestamp 1711653199
transform 1 0 340 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4478
timestamp 1711653199
transform 1 0 292 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_4479
timestamp 1711653199
transform 1 0 468 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4480
timestamp 1711653199
transform 1 0 316 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4481
timestamp 1711653199
transform 1 0 348 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4482
timestamp 1711653199
transform 1 0 260 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4483
timestamp 1711653199
transform 1 0 284 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4484
timestamp 1711653199
transform 1 0 220 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4485
timestamp 1711653199
transform 1 0 860 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4486
timestamp 1711653199
transform 1 0 564 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4487
timestamp 1711653199
transform 1 0 532 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4488
timestamp 1711653199
transform 1 0 692 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4489
timestamp 1711653199
transform 1 0 460 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4490
timestamp 1711653199
transform 1 0 188 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_4491
timestamp 1711653199
transform 1 0 108 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_4492
timestamp 1711653199
transform 1 0 180 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4493
timestamp 1711653199
transform 1 0 116 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4494
timestamp 1711653199
transform 1 0 164 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4495
timestamp 1711653199
transform 1 0 148 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4496
timestamp 1711653199
transform 1 0 132 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4497
timestamp 1711653199
transform 1 0 132 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_4498
timestamp 1711653199
transform 1 0 116 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_4499
timestamp 1711653199
transform 1 0 92 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4500
timestamp 1711653199
transform 1 0 188 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4501
timestamp 1711653199
transform 1 0 116 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4502
timestamp 1711653199
transform 1 0 148 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_4503
timestamp 1711653199
transform 1 0 116 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_4504
timestamp 1711653199
transform 1 0 132 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4505
timestamp 1711653199
transform 1 0 132 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_4506
timestamp 1711653199
transform 1 0 308 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4507
timestamp 1711653199
transform 1 0 276 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4508
timestamp 1711653199
transform 1 0 220 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4509
timestamp 1711653199
transform 1 0 116 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4510
timestamp 1711653199
transform 1 0 116 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4511
timestamp 1711653199
transform 1 0 100 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4512
timestamp 1711653199
transform 1 0 68 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4513
timestamp 1711653199
transform 1 0 108 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4514
timestamp 1711653199
transform 1 0 108 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_4515
timestamp 1711653199
transform 1 0 100 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4516
timestamp 1711653199
transform 1 0 100 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4517
timestamp 1711653199
transform 1 0 100 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4518
timestamp 1711653199
transform 1 0 100 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4519
timestamp 1711653199
transform 1 0 100 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4520
timestamp 1711653199
transform 1 0 92 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4521
timestamp 1711653199
transform 1 0 380 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4522
timestamp 1711653199
transform 1 0 84 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4523
timestamp 1711653199
transform 1 0 188 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4524
timestamp 1711653199
transform 1 0 132 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4525
timestamp 1711653199
transform 1 0 2972 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4526
timestamp 1711653199
transform 1 0 2924 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4527
timestamp 1711653199
transform 1 0 2924 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4528
timestamp 1711653199
transform 1 0 2500 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4529
timestamp 1711653199
transform 1 0 1852 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4530
timestamp 1711653199
transform 1 0 1836 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4531
timestamp 1711653199
transform 1 0 1508 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4532
timestamp 1711653199
transform 1 0 1092 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4533
timestamp 1711653199
transform 1 0 1092 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4534
timestamp 1711653199
transform 1 0 916 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_4535
timestamp 1711653199
transform 1 0 900 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4536
timestamp 1711653199
transform 1 0 900 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4537
timestamp 1711653199
transform 1 0 652 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4538
timestamp 1711653199
transform 1 0 652 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4539
timestamp 1711653199
transform 1 0 500 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4540
timestamp 1711653199
transform 1 0 284 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4541
timestamp 1711653199
transform 1 0 212 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4542
timestamp 1711653199
transform 1 0 756 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4543
timestamp 1711653199
transform 1 0 388 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4544
timestamp 1711653199
transform 1 0 2324 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4545
timestamp 1711653199
transform 1 0 2300 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4546
timestamp 1711653199
transform 1 0 2300 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4547
timestamp 1711653199
transform 1 0 2220 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4548
timestamp 1711653199
transform 1 0 2148 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4549
timestamp 1711653199
transform 1 0 2148 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4550
timestamp 1711653199
transform 1 0 2124 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4551
timestamp 1711653199
transform 1 0 2124 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4552
timestamp 1711653199
transform 1 0 1684 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4553
timestamp 1711653199
transform 1 0 1668 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4554
timestamp 1711653199
transform 1 0 1668 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_4555
timestamp 1711653199
transform 1 0 1292 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4556
timestamp 1711653199
transform 1 0 1244 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4557
timestamp 1711653199
transform 1 0 1236 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4558
timestamp 1711653199
transform 1 0 876 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4559
timestamp 1711653199
transform 1 0 124 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4560
timestamp 1711653199
transform 1 0 124 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4561
timestamp 1711653199
transform 1 0 84 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_4562
timestamp 1711653199
transform 1 0 84 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4563
timestamp 1711653199
transform 1 0 116 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4564
timestamp 1711653199
transform 1 0 92 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4565
timestamp 1711653199
transform 1 0 356 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4566
timestamp 1711653199
transform 1 0 148 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4567
timestamp 1711653199
transform 1 0 148 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4568
timestamp 1711653199
transform 1 0 84 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4569
timestamp 1711653199
transform 1 0 164 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_4570
timestamp 1711653199
transform 1 0 124 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_4571
timestamp 1711653199
transform 1 0 404 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4572
timestamp 1711653199
transform 1 0 388 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4573
timestamp 1711653199
transform 1 0 388 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4574
timestamp 1711653199
transform 1 0 356 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4575
timestamp 1711653199
transform 1 0 820 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4576
timestamp 1711653199
transform 1 0 396 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4577
timestamp 1711653199
transform 1 0 1436 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4578
timestamp 1711653199
transform 1 0 836 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4579
timestamp 1711653199
transform 1 0 836 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4580
timestamp 1711653199
transform 1 0 740 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4581
timestamp 1711653199
transform 1 0 684 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4582
timestamp 1711653199
transform 1 0 596 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4583
timestamp 1711653199
transform 1 0 532 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4584
timestamp 1711653199
transform 1 0 452 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4585
timestamp 1711653199
transform 1 0 476 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_4586
timestamp 1711653199
transform 1 0 460 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_4587
timestamp 1711653199
transform 1 0 572 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4588
timestamp 1711653199
transform 1 0 348 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_4589
timestamp 1711653199
transform 1 0 212 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4590
timestamp 1711653199
transform 1 0 132 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_4591
timestamp 1711653199
transform 1 0 228 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4592
timestamp 1711653199
transform 1 0 188 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_4593
timestamp 1711653199
transform 1 0 476 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4594
timestamp 1711653199
transform 1 0 460 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4595
timestamp 1711653199
transform 1 0 316 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4596
timestamp 1711653199
transform 1 0 156 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4597
timestamp 1711653199
transform 1 0 140 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4598
timestamp 1711653199
transform 1 0 140 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_4599
timestamp 1711653199
transform 1 0 140 0 1 1475
box -3 -3 3 3
use M3_M2  M3_M2_4600
timestamp 1711653199
transform 1 0 924 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4601
timestamp 1711653199
transform 1 0 460 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4602
timestamp 1711653199
transform 1 0 1540 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4603
timestamp 1711653199
transform 1 0 1436 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4604
timestamp 1711653199
transform 1 0 1428 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4605
timestamp 1711653199
transform 1 0 764 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4606
timestamp 1711653199
transform 1 0 764 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4607
timestamp 1711653199
transform 1 0 396 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4608
timestamp 1711653199
transform 1 0 2068 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4609
timestamp 1711653199
transform 1 0 1668 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4610
timestamp 1711653199
transform 1 0 1668 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4611
timestamp 1711653199
transform 1 0 1444 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4612
timestamp 1711653199
transform 1 0 1444 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4613
timestamp 1711653199
transform 1 0 1028 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4614
timestamp 1711653199
transform 1 0 1028 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4615
timestamp 1711653199
transform 1 0 916 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4616
timestamp 1711653199
transform 1 0 948 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4617
timestamp 1711653199
transform 1 0 884 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4618
timestamp 1711653199
transform 1 0 2404 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4619
timestamp 1711653199
transform 1 0 2388 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4620
timestamp 1711653199
transform 1 0 2084 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4621
timestamp 1711653199
transform 1 0 1740 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4622
timestamp 1711653199
transform 1 0 1700 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4623
timestamp 1711653199
transform 1 0 1268 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4624
timestamp 1711653199
transform 1 0 2116 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4625
timestamp 1711653199
transform 1 0 1964 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4626
timestamp 1711653199
transform 1 0 1044 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4627
timestamp 1711653199
transform 1 0 1044 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4628
timestamp 1711653199
transform 1 0 868 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4629
timestamp 1711653199
transform 1 0 572 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4630
timestamp 1711653199
transform 1 0 548 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4631
timestamp 1711653199
transform 1 0 484 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4632
timestamp 1711653199
transform 1 0 580 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_4633
timestamp 1711653199
transform 1 0 556 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4634
timestamp 1711653199
transform 1 0 556 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4635
timestamp 1711653199
transform 1 0 524 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4636
timestamp 1711653199
transform 1 0 748 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4637
timestamp 1711653199
transform 1 0 684 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4638
timestamp 1711653199
transform 1 0 684 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4639
timestamp 1711653199
transform 1 0 516 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4640
timestamp 1711653199
transform 1 0 620 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4641
timestamp 1711653199
transform 1 0 580 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4642
timestamp 1711653199
transform 1 0 596 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4643
timestamp 1711653199
transform 1 0 460 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4644
timestamp 1711653199
transform 1 0 1036 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4645
timestamp 1711653199
transform 1 0 876 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_4646
timestamp 1711653199
transform 1 0 876 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_4647
timestamp 1711653199
transform 1 0 564 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_4648
timestamp 1711653199
transform 1 0 524 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4649
timestamp 1711653199
transform 1 0 500 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4650
timestamp 1711653199
transform 1 0 924 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4651
timestamp 1711653199
transform 1 0 868 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4652
timestamp 1711653199
transform 1 0 868 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4653
timestamp 1711653199
transform 1 0 748 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_4654
timestamp 1711653199
transform 1 0 668 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_4655
timestamp 1711653199
transform 1 0 740 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4656
timestamp 1711653199
transform 1 0 676 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_4657
timestamp 1711653199
transform 1 0 828 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_4658
timestamp 1711653199
transform 1 0 740 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4659
timestamp 1711653199
transform 1 0 844 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4660
timestamp 1711653199
transform 1 0 724 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_4661
timestamp 1711653199
transform 1 0 908 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4662
timestamp 1711653199
transform 1 0 884 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4663
timestamp 1711653199
transform 1 0 1108 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4664
timestamp 1711653199
transform 1 0 996 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4665
timestamp 1711653199
transform 1 0 2372 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4666
timestamp 1711653199
transform 1 0 2284 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4667
timestamp 1711653199
transform 1 0 2284 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4668
timestamp 1711653199
transform 1 0 2268 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_4669
timestamp 1711653199
transform 1 0 2220 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4670
timestamp 1711653199
transform 1 0 2004 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4671
timestamp 1711653199
transform 1 0 1828 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4672
timestamp 1711653199
transform 1 0 1268 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_4673
timestamp 1711653199
transform 1 0 1252 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4674
timestamp 1711653199
transform 1 0 1220 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4675
timestamp 1711653199
transform 1 0 1180 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4676
timestamp 1711653199
transform 1 0 1180 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4677
timestamp 1711653199
transform 1 0 460 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4678
timestamp 1711653199
transform 1 0 444 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_4679
timestamp 1711653199
transform 1 0 484 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4680
timestamp 1711653199
transform 1 0 428 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4681
timestamp 1711653199
transform 1 0 516 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4682
timestamp 1711653199
transform 1 0 388 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4683
timestamp 1711653199
transform 1 0 420 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4684
timestamp 1711653199
transform 1 0 404 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4685
timestamp 1711653199
transform 1 0 852 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4686
timestamp 1711653199
transform 1 0 708 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4687
timestamp 1711653199
transform 1 0 708 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_4688
timestamp 1711653199
transform 1 0 652 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4689
timestamp 1711653199
transform 1 0 580 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4690
timestamp 1711653199
transform 1 0 580 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4691
timestamp 1711653199
transform 1 0 468 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_4692
timestamp 1711653199
transform 1 0 468 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4693
timestamp 1711653199
transform 1 0 852 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_4694
timestamp 1711653199
transform 1 0 716 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4695
timestamp 1711653199
transform 1 0 700 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4696
timestamp 1711653199
transform 1 0 700 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_4697
timestamp 1711653199
transform 1 0 700 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4698
timestamp 1711653199
transform 1 0 492 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4699
timestamp 1711653199
transform 1 0 436 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_4700
timestamp 1711653199
transform 1 0 740 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4701
timestamp 1711653199
transform 1 0 724 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4702
timestamp 1711653199
transform 1 0 684 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_4703
timestamp 1711653199
transform 1 0 540 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_4704
timestamp 1711653199
transform 1 0 596 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4705
timestamp 1711653199
transform 1 0 564 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_4706
timestamp 1711653199
transform 1 0 628 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_4707
timestamp 1711653199
transform 1 0 580 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_4708
timestamp 1711653199
transform 1 0 516 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_4709
timestamp 1711653199
transform 1 0 444 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_4710
timestamp 1711653199
transform 1 0 724 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4711
timestamp 1711653199
transform 1 0 436 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4712
timestamp 1711653199
transform 1 0 596 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_4713
timestamp 1711653199
transform 1 0 556 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_4714
timestamp 1711653199
transform 1 0 804 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4715
timestamp 1711653199
transform 1 0 716 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4716
timestamp 1711653199
transform 1 0 684 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4717
timestamp 1711653199
transform 1 0 636 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4718
timestamp 1711653199
transform 1 0 612 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4719
timestamp 1711653199
transform 1 0 612 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4720
timestamp 1711653199
transform 1 0 556 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4721
timestamp 1711653199
transform 1 0 516 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4722
timestamp 1711653199
transform 1 0 620 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4723
timestamp 1711653199
transform 1 0 500 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_4724
timestamp 1711653199
transform 1 0 700 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_4725
timestamp 1711653199
transform 1 0 524 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4726
timestamp 1711653199
transform 1 0 900 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4727
timestamp 1711653199
transform 1 0 844 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4728
timestamp 1711653199
transform 1 0 812 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_4729
timestamp 1711653199
transform 1 0 1060 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4730
timestamp 1711653199
transform 1 0 1004 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4731
timestamp 1711653199
transform 1 0 1004 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4732
timestamp 1711653199
transform 1 0 684 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4733
timestamp 1711653199
transform 1 0 636 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4734
timestamp 1711653199
transform 1 0 1764 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4735
timestamp 1711653199
transform 1 0 1068 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_4736
timestamp 1711653199
transform 1 0 1052 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4737
timestamp 1711653199
transform 1 0 988 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_4738
timestamp 1711653199
transform 1 0 772 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4739
timestamp 1711653199
transform 1 0 612 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4740
timestamp 1711653199
transform 1 0 1204 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4741
timestamp 1711653199
transform 1 0 628 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4742
timestamp 1711653199
transform 1 0 628 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4743
timestamp 1711653199
transform 1 0 532 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4744
timestamp 1711653199
transform 1 0 484 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4745
timestamp 1711653199
transform 1 0 1780 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4746
timestamp 1711653199
transform 1 0 1380 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_4747
timestamp 1711653199
transform 1 0 1332 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4748
timestamp 1711653199
transform 1 0 980 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4749
timestamp 1711653199
transform 1 0 2268 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4750
timestamp 1711653199
transform 1 0 1844 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_4751
timestamp 1711653199
transform 1 0 2100 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4752
timestamp 1711653199
transform 1 0 1852 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4753
timestamp 1711653199
transform 1 0 1780 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4754
timestamp 1711653199
transform 1 0 1764 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4755
timestamp 1711653199
transform 1 0 1748 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4756
timestamp 1711653199
transform 1 0 1732 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_4757
timestamp 1711653199
transform 1 0 1460 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_4758
timestamp 1711653199
transform 1 0 1420 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_4759
timestamp 1711653199
transform 1 0 2188 0 1 35
box -3 -3 3 3
use M3_M2  M3_M2_4760
timestamp 1711653199
transform 1 0 1756 0 1 35
box -3 -3 3 3
use M3_M2  M3_M2_4761
timestamp 1711653199
transform 1 0 1652 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_4762
timestamp 1711653199
transform 1 0 1548 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4763
timestamp 1711653199
transform 1 0 1588 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4764
timestamp 1711653199
transform 1 0 1340 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4765
timestamp 1711653199
transform 1 0 1172 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4766
timestamp 1711653199
transform 1 0 932 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4767
timestamp 1711653199
transform 1 0 1980 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4768
timestamp 1711653199
transform 1 0 1732 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4769
timestamp 1711653199
transform 1 0 1404 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4770
timestamp 1711653199
transform 1 0 1372 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4771
timestamp 1711653199
transform 1 0 1164 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4772
timestamp 1711653199
transform 1 0 1164 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4773
timestamp 1711653199
transform 1 0 964 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4774
timestamp 1711653199
transform 1 0 644 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4775
timestamp 1711653199
transform 1 0 1644 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4776
timestamp 1711653199
transform 1 0 788 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4777
timestamp 1711653199
transform 1 0 948 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4778
timestamp 1711653199
transform 1 0 900 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4779
timestamp 1711653199
transform 1 0 876 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4780
timestamp 1711653199
transform 1 0 804 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_4781
timestamp 1711653199
transform 1 0 844 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4782
timestamp 1711653199
transform 1 0 804 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_4783
timestamp 1711653199
transform 1 0 828 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_4784
timestamp 1711653199
transform 1 0 772 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_4785
timestamp 1711653199
transform 1 0 932 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4786
timestamp 1711653199
transform 1 0 860 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4787
timestamp 1711653199
transform 1 0 852 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4788
timestamp 1711653199
transform 1 0 804 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4789
timestamp 1711653199
transform 1 0 796 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4790
timestamp 1711653199
transform 1 0 764 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_4791
timestamp 1711653199
transform 1 0 1556 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4792
timestamp 1711653199
transform 1 0 836 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_4793
timestamp 1711653199
transform 1 0 788 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4794
timestamp 1711653199
transform 1 0 516 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_4795
timestamp 1711653199
transform 1 0 868 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4796
timestamp 1711653199
transform 1 0 796 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4797
timestamp 1711653199
transform 1 0 844 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4798
timestamp 1711653199
transform 1 0 804 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_4799
timestamp 1711653199
transform 1 0 868 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4800
timestamp 1711653199
transform 1 0 748 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4801
timestamp 1711653199
transform 1 0 804 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4802
timestamp 1711653199
transform 1 0 788 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4803
timestamp 1711653199
transform 1 0 652 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4804
timestamp 1711653199
transform 1 0 596 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_4805
timestamp 1711653199
transform 1 0 596 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_4806
timestamp 1711653199
transform 1 0 500 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_4807
timestamp 1711653199
transform 1 0 452 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4808
timestamp 1711653199
transform 1 0 452 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4809
timestamp 1711653199
transform 1 0 436 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4810
timestamp 1711653199
transform 1 0 436 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_4811
timestamp 1711653199
transform 1 0 396 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4812
timestamp 1711653199
transform 1 0 396 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_4813
timestamp 1711653199
transform 1 0 388 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4814
timestamp 1711653199
transform 1 0 364 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4815
timestamp 1711653199
transform 1 0 420 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4816
timestamp 1711653199
transform 1 0 380 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_4817
timestamp 1711653199
transform 1 0 500 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_4818
timestamp 1711653199
transform 1 0 428 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4819
timestamp 1711653199
transform 1 0 388 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_4820
timestamp 1711653199
transform 1 0 444 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4821
timestamp 1711653199
transform 1 0 412 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4822
timestamp 1711653199
transform 1 0 436 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4823
timestamp 1711653199
transform 1 0 380 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_4824
timestamp 1711653199
transform 1 0 436 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4825
timestamp 1711653199
transform 1 0 412 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4826
timestamp 1711653199
transform 1 0 412 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4827
timestamp 1711653199
transform 1 0 412 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_4828
timestamp 1711653199
transform 1 0 388 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4829
timestamp 1711653199
transform 1 0 364 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_4830
timestamp 1711653199
transform 1 0 404 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4831
timestamp 1711653199
transform 1 0 380 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4832
timestamp 1711653199
transform 1 0 284 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4833
timestamp 1711653199
transform 1 0 212 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_4834
timestamp 1711653199
transform 1 0 508 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4835
timestamp 1711653199
transform 1 0 508 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4836
timestamp 1711653199
transform 1 0 468 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_4837
timestamp 1711653199
transform 1 0 468 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4838
timestamp 1711653199
transform 1 0 548 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4839
timestamp 1711653199
transform 1 0 484 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4840
timestamp 1711653199
transform 1 0 516 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4841
timestamp 1711653199
transform 1 0 476 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_4842
timestamp 1711653199
transform 1 0 812 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4843
timestamp 1711653199
transform 1 0 716 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_4844
timestamp 1711653199
transform 1 0 668 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4845
timestamp 1711653199
transform 1 0 564 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4846
timestamp 1711653199
transform 1 0 580 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4847
timestamp 1711653199
transform 1 0 276 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4848
timestamp 1711653199
transform 1 0 260 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4849
timestamp 1711653199
transform 1 0 196 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_4850
timestamp 1711653199
transform 1 0 124 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4851
timestamp 1711653199
transform 1 0 84 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_4852
timestamp 1711653199
transform 1 0 228 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4853
timestamp 1711653199
transform 1 0 148 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_4854
timestamp 1711653199
transform 1 0 308 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4855
timestamp 1711653199
transform 1 0 228 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_4856
timestamp 1711653199
transform 1 0 252 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4857
timestamp 1711653199
transform 1 0 220 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_4858
timestamp 1711653199
transform 1 0 380 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_4859
timestamp 1711653199
transform 1 0 292 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_4860
timestamp 1711653199
transform 1 0 260 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_4861
timestamp 1711653199
transform 1 0 196 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4862
timestamp 1711653199
transform 1 0 148 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_4863
timestamp 1711653199
transform 1 0 340 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4864
timestamp 1711653199
transform 1 0 284 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4865
timestamp 1711653199
transform 1 0 364 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4866
timestamp 1711653199
transform 1 0 340 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_4867
timestamp 1711653199
transform 1 0 372 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_4868
timestamp 1711653199
transform 1 0 372 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4869
timestamp 1711653199
transform 1 0 348 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4870
timestamp 1711653199
transform 1 0 340 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_4871
timestamp 1711653199
transform 1 0 324 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_4872
timestamp 1711653199
transform 1 0 316 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4873
timestamp 1711653199
transform 1 0 1332 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_4874
timestamp 1711653199
transform 1 0 300 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_4875
timestamp 1711653199
transform 1 0 196 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_4876
timestamp 1711653199
transform 1 0 3004 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_4877
timestamp 1711653199
transform 1 0 1380 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_4878
timestamp 1711653199
transform 1 0 284 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4879
timestamp 1711653199
transform 1 0 244 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4880
timestamp 1711653199
transform 1 0 244 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4881
timestamp 1711653199
transform 1 0 244 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4882
timestamp 1711653199
transform 1 0 220 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_4883
timestamp 1711653199
transform 1 0 212 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_4884
timestamp 1711653199
transform 1 0 116 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_4885
timestamp 1711653199
transform 1 0 116 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4886
timestamp 1711653199
transform 1 0 116 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_4887
timestamp 1711653199
transform 1 0 116 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_4888
timestamp 1711653199
transform 1 0 68 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4889
timestamp 1711653199
transform 1 0 68 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_4890
timestamp 1711653199
transform 1 0 380 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4891
timestamp 1711653199
transform 1 0 260 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4892
timestamp 1711653199
transform 1 0 1036 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4893
timestamp 1711653199
transform 1 0 692 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4894
timestamp 1711653199
transform 1 0 692 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4895
timestamp 1711653199
transform 1 0 596 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4896
timestamp 1711653199
transform 1 0 668 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4897
timestamp 1711653199
transform 1 0 388 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4898
timestamp 1711653199
transform 1 0 1452 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4899
timestamp 1711653199
transform 1 0 1444 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4900
timestamp 1711653199
transform 1 0 1396 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4901
timestamp 1711653199
transform 1 0 1396 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4902
timestamp 1711653199
transform 1 0 1412 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4903
timestamp 1711653199
transform 1 0 1348 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4904
timestamp 1711653199
transform 1 0 1388 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4905
timestamp 1711653199
transform 1 0 1364 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_4906
timestamp 1711653199
transform 1 0 1396 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4907
timestamp 1711653199
transform 1 0 1276 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_4908
timestamp 1711653199
transform 1 0 1276 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4909
timestamp 1711653199
transform 1 0 1252 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_4910
timestamp 1711653199
transform 1 0 2388 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4911
timestamp 1711653199
transform 1 0 2300 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4912
timestamp 1711653199
transform 1 0 2204 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4913
timestamp 1711653199
transform 1 0 1404 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4914
timestamp 1711653199
transform 1 0 1404 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4915
timestamp 1711653199
transform 1 0 1340 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4916
timestamp 1711653199
transform 1 0 1396 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4917
timestamp 1711653199
transform 1 0 1380 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_4918
timestamp 1711653199
transform 1 0 1404 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_4919
timestamp 1711653199
transform 1 0 1340 0 1 85
box -3 -3 3 3
use M3_M2  M3_M2_4920
timestamp 1711653199
transform 1 0 1476 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_4921
timestamp 1711653199
transform 1 0 1476 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_4922
timestamp 1711653199
transform 1 0 1476 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4923
timestamp 1711653199
transform 1 0 1380 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4924
timestamp 1711653199
transform 1 0 1316 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_4925
timestamp 1711653199
transform 1 0 1316 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4926
timestamp 1711653199
transform 1 0 1252 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4927
timestamp 1711653199
transform 1 0 1164 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_4928
timestamp 1711653199
transform 1 0 1476 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4929
timestamp 1711653199
transform 1 0 1444 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_4930
timestamp 1711653199
transform 1 0 2476 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4931
timestamp 1711653199
transform 1 0 2396 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4932
timestamp 1711653199
transform 1 0 2228 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_4933
timestamp 1711653199
transform 1 0 2228 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4934
timestamp 1711653199
transform 1 0 1500 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4935
timestamp 1711653199
transform 1 0 1500 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_4936
timestamp 1711653199
transform 1 0 1460 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_4937
timestamp 1711653199
transform 1 0 1388 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4938
timestamp 1711653199
transform 1 0 1188 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4939
timestamp 1711653199
transform 1 0 2012 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4940
timestamp 1711653199
transform 1 0 1516 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4941
timestamp 1711653199
transform 1 0 1476 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4942
timestamp 1711653199
transform 1 0 1268 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4943
timestamp 1711653199
transform 1 0 1332 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4944
timestamp 1711653199
transform 1 0 1180 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_4945
timestamp 1711653199
transform 1 0 1052 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4946
timestamp 1711653199
transform 1 0 964 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_4947
timestamp 1711653199
transform 1 0 1356 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4948
timestamp 1711653199
transform 1 0 1340 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4949
timestamp 1711653199
transform 1 0 1332 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_4950
timestamp 1711653199
transform 1 0 1252 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4951
timestamp 1711653199
transform 1 0 1180 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_4952
timestamp 1711653199
transform 1 0 1228 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4953
timestamp 1711653199
transform 1 0 1220 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4954
timestamp 1711653199
transform 1 0 1172 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_4955
timestamp 1711653199
transform 1 0 1124 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4956
timestamp 1711653199
transform 1 0 1100 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4957
timestamp 1711653199
transform 1 0 1100 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4958
timestamp 1711653199
transform 1 0 1044 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4959
timestamp 1711653199
transform 1 0 1044 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4960
timestamp 1711653199
transform 1 0 1044 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_4961
timestamp 1711653199
transform 1 0 996 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_4962
timestamp 1711653199
transform 1 0 996 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_4963
timestamp 1711653199
transform 1 0 1252 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4964
timestamp 1711653199
transform 1 0 1124 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_4965
timestamp 1711653199
transform 1 0 1084 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4966
timestamp 1711653199
transform 1 0 996 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_4967
timestamp 1711653199
transform 1 0 1212 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4968
timestamp 1711653199
transform 1 0 1148 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_4969
timestamp 1711653199
transform 1 0 1332 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4970
timestamp 1711653199
transform 1 0 1276 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4971
timestamp 1711653199
transform 1 0 1316 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4972
timestamp 1711653199
transform 1 0 1276 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4973
timestamp 1711653199
transform 1 0 1860 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4974
timestamp 1711653199
transform 1 0 1524 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4975
timestamp 1711653199
transform 1 0 1956 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4976
timestamp 1711653199
transform 1 0 1860 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_4977
timestamp 1711653199
transform 1 0 2892 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4978
timestamp 1711653199
transform 1 0 2860 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4979
timestamp 1711653199
transform 1 0 2764 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4980
timestamp 1711653199
transform 1 0 2668 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4981
timestamp 1711653199
transform 1 0 2668 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4982
timestamp 1711653199
transform 1 0 2612 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4983
timestamp 1711653199
transform 1 0 2324 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4984
timestamp 1711653199
transform 1 0 2148 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4985
timestamp 1711653199
transform 1 0 2148 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4986
timestamp 1711653199
transform 1 0 1948 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4987
timestamp 1711653199
transform 1 0 1652 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4988
timestamp 1711653199
transform 1 0 1572 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4989
timestamp 1711653199
transform 1 0 1572 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4990
timestamp 1711653199
transform 1 0 1564 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_4991
timestamp 1711653199
transform 1 0 1556 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4992
timestamp 1711653199
transform 1 0 1532 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_4993
timestamp 1711653199
transform 1 0 1516 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_4994
timestamp 1711653199
transform 1 0 1372 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_4995
timestamp 1711653199
transform 1 0 1332 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4996
timestamp 1711653199
transform 1 0 1276 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_4997
timestamp 1711653199
transform 1 0 1276 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4998
timestamp 1711653199
transform 1 0 1236 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_4999
timestamp 1711653199
transform 1 0 1244 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5000
timestamp 1711653199
transform 1 0 1212 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5001
timestamp 1711653199
transform 1 0 1116 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5002
timestamp 1711653199
transform 1 0 1212 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5003
timestamp 1711653199
transform 1 0 1212 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5004
timestamp 1711653199
transform 1 0 1132 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5005
timestamp 1711653199
transform 1 0 1132 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5006
timestamp 1711653199
transform 1 0 1220 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5007
timestamp 1711653199
transform 1 0 1140 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5008
timestamp 1711653199
transform 1 0 2996 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5009
timestamp 1711653199
transform 1 0 2972 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5010
timestamp 1711653199
transform 1 0 2972 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5011
timestamp 1711653199
transform 1 0 2860 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5012
timestamp 1711653199
transform 1 0 2420 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5013
timestamp 1711653199
transform 1 0 2372 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5014
timestamp 1711653199
transform 1 0 2372 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5015
timestamp 1711653199
transform 1 0 2260 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5016
timestamp 1711653199
transform 1 0 2260 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5017
timestamp 1711653199
transform 1 0 2180 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5018
timestamp 1711653199
transform 1 0 1428 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5019
timestamp 1711653199
transform 1 0 1764 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_5020
timestamp 1711653199
transform 1 0 1700 0 1 2075
box -3 -3 3 3
use M3_M2  M3_M2_5021
timestamp 1711653199
transform 1 0 2380 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5022
timestamp 1711653199
transform 1 0 2116 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_5023
timestamp 1711653199
transform 1 0 2068 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5024
timestamp 1711653199
transform 1 0 2068 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_5025
timestamp 1711653199
transform 1 0 1732 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5026
timestamp 1711653199
transform 1 0 1412 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5027
timestamp 1711653199
transform 1 0 1116 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5028
timestamp 1711653199
transform 1 0 1076 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_5029
timestamp 1711653199
transform 1 0 1076 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_5030
timestamp 1711653199
transform 1 0 1012 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_5031
timestamp 1711653199
transform 1 0 1004 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_5032
timestamp 1711653199
transform 1 0 1068 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5033
timestamp 1711653199
transform 1 0 1052 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_5034
timestamp 1711653199
transform 1 0 1156 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5035
timestamp 1711653199
transform 1 0 1132 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5036
timestamp 1711653199
transform 1 0 1116 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5037
timestamp 1711653199
transform 1 0 1020 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5038
timestamp 1711653199
transform 1 0 1164 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5039
timestamp 1711653199
transform 1 0 1124 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_5040
timestamp 1711653199
transform 1 0 1100 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5041
timestamp 1711653199
transform 1 0 1068 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_5042
timestamp 1711653199
transform 1 0 1060 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5043
timestamp 1711653199
transform 1 0 980 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_5044
timestamp 1711653199
transform 1 0 1940 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_5045
timestamp 1711653199
transform 1 0 1628 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_5046
timestamp 1711653199
transform 1 0 1612 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_5047
timestamp 1711653199
transform 1 0 1092 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_5048
timestamp 1711653199
transform 1 0 1180 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5049
timestamp 1711653199
transform 1 0 1164 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5050
timestamp 1711653199
transform 1 0 1044 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5051
timestamp 1711653199
transform 1 0 964 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_5052
timestamp 1711653199
transform 1 0 1116 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5053
timestamp 1711653199
transform 1 0 1068 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_5054
timestamp 1711653199
transform 1 0 2468 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5055
timestamp 1711653199
transform 1 0 2356 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5056
timestamp 1711653199
transform 1 0 2092 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5057
timestamp 1711653199
transform 1 0 1348 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5058
timestamp 1711653199
transform 1 0 1844 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5059
timestamp 1711653199
transform 1 0 1780 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5060
timestamp 1711653199
transform 1 0 2148 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5061
timestamp 1711653199
transform 1 0 2044 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5062
timestamp 1711653199
transform 1 0 1812 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5063
timestamp 1711653199
transform 1 0 2428 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_5064
timestamp 1711653199
transform 1 0 2268 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_5065
timestamp 1711653199
transform 1 0 2532 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_5066
timestamp 1711653199
transform 1 0 2412 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_5067
timestamp 1711653199
transform 1 0 2564 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_5068
timestamp 1711653199
transform 1 0 2500 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_5069
timestamp 1711653199
transform 1 0 2252 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_5070
timestamp 1711653199
transform 1 0 2052 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5071
timestamp 1711653199
transform 1 0 2052 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_5072
timestamp 1711653199
transform 1 0 2036 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5073
timestamp 1711653199
transform 1 0 1972 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_5074
timestamp 1711653199
transform 1 0 2604 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5075
timestamp 1711653199
transform 1 0 2540 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5076
timestamp 1711653199
transform 1 0 2564 0 1 65
box -3 -3 3 3
use M3_M2  M3_M2_5077
timestamp 1711653199
transform 1 0 2244 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_5078
timestamp 1711653199
transform 1 0 2532 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5079
timestamp 1711653199
transform 1 0 2436 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5080
timestamp 1711653199
transform 1 0 2380 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_5081
timestamp 1711653199
transform 1 0 2132 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_5082
timestamp 1711653199
transform 1 0 2348 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_5083
timestamp 1711653199
transform 1 0 2300 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_5084
timestamp 1711653199
transform 1 0 2220 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5085
timestamp 1711653199
transform 1 0 2196 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5086
timestamp 1711653199
transform 1 0 2684 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5087
timestamp 1711653199
transform 1 0 2636 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5088
timestamp 1711653199
transform 1 0 2548 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5089
timestamp 1711653199
transform 1 0 2548 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_5090
timestamp 1711653199
transform 1 0 2540 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_5091
timestamp 1711653199
transform 1 0 2516 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5092
timestamp 1711653199
transform 1 0 2484 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_5093
timestamp 1711653199
transform 1 0 2484 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5094
timestamp 1711653199
transform 1 0 2268 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5095
timestamp 1711653199
transform 1 0 2252 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5096
timestamp 1711653199
transform 1 0 2012 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5097
timestamp 1711653199
transform 1 0 2772 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5098
timestamp 1711653199
transform 1 0 2684 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5099
timestamp 1711653199
transform 1 0 2580 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5100
timestamp 1711653199
transform 1 0 2580 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5101
timestamp 1711653199
transform 1 0 2292 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5102
timestamp 1711653199
transform 1 0 2004 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5103
timestamp 1711653199
transform 1 0 1596 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5104
timestamp 1711653199
transform 1 0 1980 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5105
timestamp 1711653199
transform 1 0 1932 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_5106
timestamp 1711653199
transform 1 0 3220 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5107
timestamp 1711653199
transform 1 0 3220 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_5108
timestamp 1711653199
transform 1 0 3180 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5109
timestamp 1711653199
transform 1 0 3172 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5110
timestamp 1711653199
transform 1 0 3116 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_5111
timestamp 1711653199
transform 1 0 2316 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_5112
timestamp 1711653199
transform 1 0 3196 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5113
timestamp 1711653199
transform 1 0 3052 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_5114
timestamp 1711653199
transform 1 0 3188 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5115
timestamp 1711653199
transform 1 0 3148 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5116
timestamp 1711653199
transform 1 0 3172 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_5117
timestamp 1711653199
transform 1 0 3132 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_5118
timestamp 1711653199
transform 1 0 3172 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_5119
timestamp 1711653199
transform 1 0 3060 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5120
timestamp 1711653199
transform 1 0 3044 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5121
timestamp 1711653199
transform 1 0 3044 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_5122
timestamp 1711653199
transform 1 0 2956 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5123
timestamp 1711653199
transform 1 0 2956 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_5124
timestamp 1711653199
transform 1 0 2556 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5125
timestamp 1711653199
transform 1 0 3204 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5126
timestamp 1711653199
transform 1 0 3132 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_5127
timestamp 1711653199
transform 1 0 3092 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_5128
timestamp 1711653199
transform 1 0 3068 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_5129
timestamp 1711653199
transform 1 0 3108 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5130
timestamp 1711653199
transform 1 0 3036 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5131
timestamp 1711653199
transform 1 0 3052 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5132
timestamp 1711653199
transform 1 0 2980 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5133
timestamp 1711653199
transform 1 0 3124 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5134
timestamp 1711653199
transform 1 0 3076 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5135
timestamp 1711653199
transform 1 0 3060 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5136
timestamp 1711653199
transform 1 0 3004 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_5137
timestamp 1711653199
transform 1 0 3004 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_5138
timestamp 1711653199
transform 1 0 2948 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_5139
timestamp 1711653199
transform 1 0 3124 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5140
timestamp 1711653199
transform 1 0 3076 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5141
timestamp 1711653199
transform 1 0 3132 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_5142
timestamp 1711653199
transform 1 0 3044 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_5143
timestamp 1711653199
transform 1 0 3148 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5144
timestamp 1711653199
transform 1 0 2548 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5145
timestamp 1711653199
transform 1 0 2548 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5146
timestamp 1711653199
transform 1 0 2460 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5147
timestamp 1711653199
transform 1 0 3396 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_5148
timestamp 1711653199
transform 1 0 3396 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5149
timestamp 1711653199
transform 1 0 3396 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_5150
timestamp 1711653199
transform 1 0 3380 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5151
timestamp 1711653199
transform 1 0 3300 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_5152
timestamp 1711653199
transform 1 0 3084 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_5153
timestamp 1711653199
transform 1 0 3084 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5154
timestamp 1711653199
transform 1 0 2620 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_5155
timestamp 1711653199
transform 1 0 3396 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_5156
timestamp 1711653199
transform 1 0 3284 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_5157
timestamp 1711653199
transform 1 0 3340 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5158
timestamp 1711653199
transform 1 0 3324 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5159
timestamp 1711653199
transform 1 0 3284 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_5160
timestamp 1711653199
transform 1 0 3228 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_5161
timestamp 1711653199
transform 1 0 3324 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5162
timestamp 1711653199
transform 1 0 3276 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_5163
timestamp 1711653199
transform 1 0 3228 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5164
timestamp 1711653199
transform 1 0 3228 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5165
timestamp 1711653199
transform 1 0 3292 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_5166
timestamp 1711653199
transform 1 0 3220 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_5167
timestamp 1711653199
transform 1 0 3308 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5168
timestamp 1711653199
transform 1 0 3252 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5169
timestamp 1711653199
transform 1 0 3196 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5170
timestamp 1711653199
transform 1 0 3188 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5171
timestamp 1711653199
transform 1 0 3172 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_5172
timestamp 1711653199
transform 1 0 3172 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5173
timestamp 1711653199
transform 1 0 3132 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_5174
timestamp 1711653199
transform 1 0 3132 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_5175
timestamp 1711653199
transform 1 0 3188 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5176
timestamp 1711653199
transform 1 0 3172 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5177
timestamp 1711653199
transform 1 0 3172 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5178
timestamp 1711653199
transform 1 0 3148 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5179
timestamp 1711653199
transform 1 0 3268 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5180
timestamp 1711653199
transform 1 0 3196 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5181
timestamp 1711653199
transform 1 0 2988 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5182
timestamp 1711653199
transform 1 0 2988 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5183
timestamp 1711653199
transform 1 0 2932 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5184
timestamp 1711653199
transform 1 0 2932 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5185
timestamp 1711653199
transform 1 0 2820 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5186
timestamp 1711653199
transform 1 0 2812 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5187
timestamp 1711653199
transform 1 0 2572 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5188
timestamp 1711653199
transform 1 0 2564 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_5189
timestamp 1711653199
transform 1 0 2380 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5190
timestamp 1711653199
transform 1 0 3164 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5191
timestamp 1711653199
transform 1 0 3020 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5192
timestamp 1711653199
transform 1 0 3020 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_5193
timestamp 1711653199
transform 1 0 2852 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5194
timestamp 1711653199
transform 1 0 2852 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_5195
timestamp 1711653199
transform 1 0 2372 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5196
timestamp 1711653199
transform 1 0 3372 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_5197
timestamp 1711653199
transform 1 0 3348 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5198
timestamp 1711653199
transform 1 0 3268 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5199
timestamp 1711653199
transform 1 0 3268 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_5200
timestamp 1711653199
transform 1 0 3172 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_5201
timestamp 1711653199
transform 1 0 2676 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_5202
timestamp 1711653199
transform 1 0 3212 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5203
timestamp 1711653199
transform 1 0 3156 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_5204
timestamp 1711653199
transform 1 0 3148 0 1 804
box -3 -3 3 3
use M3_M2  M3_M2_5205
timestamp 1711653199
transform 1 0 3148 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_5206
timestamp 1711653199
transform 1 0 3228 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_5207
timestamp 1711653199
transform 1 0 3156 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_5208
timestamp 1711653199
transform 1 0 3380 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_5209
timestamp 1711653199
transform 1 0 3356 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5210
timestamp 1711653199
transform 1 0 3348 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_5211
timestamp 1711653199
transform 1 0 3348 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_5212
timestamp 1711653199
transform 1 0 3340 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_5213
timestamp 1711653199
transform 1 0 3340 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_5214
timestamp 1711653199
transform 1 0 3396 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5215
timestamp 1711653199
transform 1 0 3340 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5216
timestamp 1711653199
transform 1 0 3380 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5217
timestamp 1711653199
transform 1 0 3380 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5218
timestamp 1711653199
transform 1 0 3340 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_5219
timestamp 1711653199
transform 1 0 3252 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_5220
timestamp 1711653199
transform 1 0 3236 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_5221
timestamp 1711653199
transform 1 0 3164 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_5222
timestamp 1711653199
transform 1 0 2876 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_5223
timestamp 1711653199
transform 1 0 3316 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5224
timestamp 1711653199
transform 1 0 3252 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_5225
timestamp 1711653199
transform 1 0 3268 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5226
timestamp 1711653199
transform 1 0 3196 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_5227
timestamp 1711653199
transform 1 0 3372 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_5228
timestamp 1711653199
transform 1 0 3372 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_5229
timestamp 1711653199
transform 1 0 3356 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5230
timestamp 1711653199
transform 1 0 3132 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5231
timestamp 1711653199
transform 1 0 3396 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5232
timestamp 1711653199
transform 1 0 3348 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5233
timestamp 1711653199
transform 1 0 2820 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5234
timestamp 1711653199
transform 1 0 2724 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5235
timestamp 1711653199
transform 1 0 2708 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5236
timestamp 1711653199
transform 1 0 2700 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5237
timestamp 1711653199
transform 1 0 2508 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5238
timestamp 1711653199
transform 1 0 3140 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5239
timestamp 1711653199
transform 1 0 2836 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5240
timestamp 1711653199
transform 1 0 3388 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5241
timestamp 1711653199
transform 1 0 3388 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_5242
timestamp 1711653199
transform 1 0 2772 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_5243
timestamp 1711653199
transform 1 0 2436 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5244
timestamp 1711653199
transform 1 0 2764 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_5245
timestamp 1711653199
transform 1 0 2708 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_5246
timestamp 1711653199
transform 1 0 2700 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_5247
timestamp 1711653199
transform 1 0 2628 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_5248
timestamp 1711653199
transform 1 0 2868 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_5249
timestamp 1711653199
transform 1 0 2836 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_5250
timestamp 1711653199
transform 1 0 2796 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_5251
timestamp 1711653199
transform 1 0 2772 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_5252
timestamp 1711653199
transform 1 0 2764 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_5253
timestamp 1711653199
transform 1 0 2908 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_5254
timestamp 1711653199
transform 1 0 2860 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_5255
timestamp 1711653199
transform 1 0 2756 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_5256
timestamp 1711653199
transform 1 0 2636 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_5257
timestamp 1711653199
transform 1 0 2756 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5258
timestamp 1711653199
transform 1 0 2692 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5259
timestamp 1711653199
transform 1 0 2692 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5260
timestamp 1711653199
transform 1 0 2620 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5261
timestamp 1711653199
transform 1 0 2980 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_5262
timestamp 1711653199
transform 1 0 2940 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_5263
timestamp 1711653199
transform 1 0 2860 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_5264
timestamp 1711653199
transform 1 0 2724 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_5265
timestamp 1711653199
transform 1 0 3028 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5266
timestamp 1711653199
transform 1 0 3028 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5267
timestamp 1711653199
transform 1 0 3004 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5268
timestamp 1711653199
transform 1 0 2892 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5269
timestamp 1711653199
transform 1 0 2892 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5270
timestamp 1711653199
transform 1 0 2884 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5271
timestamp 1711653199
transform 1 0 2788 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5272
timestamp 1711653199
transform 1 0 2708 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5273
timestamp 1711653199
transform 1 0 2708 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5274
timestamp 1711653199
transform 1 0 2644 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5275
timestamp 1711653199
transform 1 0 2644 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_5276
timestamp 1711653199
transform 1 0 2636 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_5277
timestamp 1711653199
transform 1 0 2476 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5278
timestamp 1711653199
transform 1 0 2820 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_5279
timestamp 1711653199
transform 1 0 2748 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_5280
timestamp 1711653199
transform 1 0 3156 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5281
timestamp 1711653199
transform 1 0 2988 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_5282
timestamp 1711653199
transform 1 0 3148 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5283
timestamp 1711653199
transform 1 0 3004 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_5284
timestamp 1711653199
transform 1 0 2852 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_5285
timestamp 1711653199
transform 1 0 2828 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5286
timestamp 1711653199
transform 1 0 2828 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_5287
timestamp 1711653199
transform 1 0 2788 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5288
timestamp 1711653199
transform 1 0 2780 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5289
timestamp 1711653199
transform 1 0 2852 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_5290
timestamp 1711653199
transform 1 0 2692 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5291
timestamp 1711653199
transform 1 0 2652 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_5292
timestamp 1711653199
transform 1 0 2652 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_5293
timestamp 1711653199
transform 1 0 3228 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_5294
timestamp 1711653199
transform 1 0 2916 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_5295
timestamp 1711653199
transform 1 0 2916 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_5296
timestamp 1711653199
transform 1 0 2908 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5297
timestamp 1711653199
transform 1 0 2844 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5298
timestamp 1711653199
transform 1 0 2844 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_5299
timestamp 1711653199
transform 1 0 2732 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_5300
timestamp 1711653199
transform 1 0 2804 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5301
timestamp 1711653199
transform 1 0 2740 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5302
timestamp 1711653199
transform 1 0 2708 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5303
timestamp 1711653199
transform 1 0 2444 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5304
timestamp 1711653199
transform 1 0 2956 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5305
timestamp 1711653199
transform 1 0 2892 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5306
timestamp 1711653199
transform 1 0 2892 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5307
timestamp 1711653199
transform 1 0 2684 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5308
timestamp 1711653199
transform 1 0 2684 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5309
timestamp 1711653199
transform 1 0 2548 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5310
timestamp 1711653199
transform 1 0 2340 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5311
timestamp 1711653199
transform 1 0 2484 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5312
timestamp 1711653199
transform 1 0 2436 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5313
timestamp 1711653199
transform 1 0 2412 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5314
timestamp 1711653199
transform 1 0 2812 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5315
timestamp 1711653199
transform 1 0 2788 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5316
timestamp 1711653199
transform 1 0 2812 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_5317
timestamp 1711653199
transform 1 0 2748 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_5318
timestamp 1711653199
transform 1 0 2740 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5319
timestamp 1711653199
transform 1 0 2684 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_5320
timestamp 1711653199
transform 1 0 2684 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5321
timestamp 1711653199
transform 1 0 2348 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_5322
timestamp 1711653199
transform 1 0 2716 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5323
timestamp 1711653199
transform 1 0 2700 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5324
timestamp 1711653199
transform 1 0 2772 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_5325
timestamp 1711653199
transform 1 0 2732 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_5326
timestamp 1711653199
transform 1 0 2780 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5327
timestamp 1711653199
transform 1 0 2748 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5328
timestamp 1711653199
transform 1 0 2772 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5329
timestamp 1711653199
transform 1 0 2700 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5330
timestamp 1711653199
transform 1 0 2732 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_5331
timestamp 1711653199
transform 1 0 2676 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_5332
timestamp 1711653199
transform 1 0 2668 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5333
timestamp 1711653199
transform 1 0 2628 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_5334
timestamp 1711653199
transform 1 0 2628 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_5335
timestamp 1711653199
transform 1 0 2516 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5336
timestamp 1711653199
transform 1 0 2740 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_5337
timestamp 1711653199
transform 1 0 2716 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_5338
timestamp 1711653199
transform 1 0 2716 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5339
timestamp 1711653199
transform 1 0 2692 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5340
timestamp 1711653199
transform 1 0 2668 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5341
timestamp 1711653199
transform 1 0 2612 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5342
timestamp 1711653199
transform 1 0 2732 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5343
timestamp 1711653199
transform 1 0 2596 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5344
timestamp 1711653199
transform 1 0 2700 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_5345
timestamp 1711653199
transform 1 0 2564 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_5346
timestamp 1711653199
transform 1 0 2692 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5347
timestamp 1711653199
transform 1 0 2644 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5348
timestamp 1711653199
transform 1 0 2652 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5349
timestamp 1711653199
transform 1 0 2452 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5350
timestamp 1711653199
transform 1 0 2356 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5351
timestamp 1711653199
transform 1 0 2348 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5352
timestamp 1711653199
transform 1 0 2324 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5353
timestamp 1711653199
transform 1 0 2324 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5354
timestamp 1711653199
transform 1 0 3012 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5355
timestamp 1711653199
transform 1 0 2820 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5356
timestamp 1711653199
transform 1 0 2652 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5357
timestamp 1711653199
transform 1 0 2692 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5358
timestamp 1711653199
transform 1 0 2620 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5359
timestamp 1711653199
transform 1 0 2812 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5360
timestamp 1711653199
transform 1 0 2628 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5361
timestamp 1711653199
transform 1 0 2644 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5362
timestamp 1711653199
transform 1 0 2564 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5363
timestamp 1711653199
transform 1 0 2588 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5364
timestamp 1711653199
transform 1 0 2348 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5365
timestamp 1711653199
transform 1 0 2468 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5366
timestamp 1711653199
transform 1 0 2396 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_5367
timestamp 1711653199
transform 1 0 2660 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5368
timestamp 1711653199
transform 1 0 2460 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5369
timestamp 1711653199
transform 1 0 2940 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5370
timestamp 1711653199
transform 1 0 2460 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5371
timestamp 1711653199
transform 1 0 2940 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5372
timestamp 1711653199
transform 1 0 2900 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5373
timestamp 1711653199
transform 1 0 2812 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5374
timestamp 1711653199
transform 1 0 2716 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_5375
timestamp 1711653199
transform 1 0 2940 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5376
timestamp 1711653199
transform 1 0 2844 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_5377
timestamp 1711653199
transform 1 0 2924 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5378
timestamp 1711653199
transform 1 0 2820 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_5379
timestamp 1711653199
transform 1 0 2956 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_5380
timestamp 1711653199
transform 1 0 2868 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_5381
timestamp 1711653199
transform 1 0 2812 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_5382
timestamp 1711653199
transform 1 0 3108 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_5383
timestamp 1711653199
transform 1 0 2972 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_5384
timestamp 1711653199
transform 1 0 2924 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_5385
timestamp 1711653199
transform 1 0 2884 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_5386
timestamp 1711653199
transform 1 0 2884 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_5387
timestamp 1711653199
transform 1 0 2692 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5388
timestamp 1711653199
transform 1 0 2644 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5389
timestamp 1711653199
transform 1 0 2684 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5390
timestamp 1711653199
transform 1 0 2564 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5391
timestamp 1711653199
transform 1 0 2596 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5392
timestamp 1711653199
transform 1 0 2532 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5393
timestamp 1711653199
transform 1 0 2572 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5394
timestamp 1711653199
transform 1 0 2508 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5395
timestamp 1711653199
transform 1 0 2644 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5396
timestamp 1711653199
transform 1 0 2572 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_5397
timestamp 1711653199
transform 1 0 2596 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_5398
timestamp 1711653199
transform 1 0 2524 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_5399
timestamp 1711653199
transform 1 0 2644 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5400
timestamp 1711653199
transform 1 0 2556 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_5401
timestamp 1711653199
transform 1 0 2708 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5402
timestamp 1711653199
transform 1 0 2708 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5403
timestamp 1711653199
transform 1 0 2668 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5404
timestamp 1711653199
transform 1 0 2660 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5405
timestamp 1711653199
transform 1 0 2580 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5406
timestamp 1711653199
transform 1 0 2444 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5407
timestamp 1711653199
transform 1 0 2660 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5408
timestamp 1711653199
transform 1 0 2588 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5409
timestamp 1711653199
transform 1 0 2660 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5410
timestamp 1711653199
transform 1 0 2540 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5411
timestamp 1711653199
transform 1 0 2556 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5412
timestamp 1711653199
transform 1 0 2460 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5413
timestamp 1711653199
transform 1 0 2916 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5414
timestamp 1711653199
transform 1 0 2900 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_5415
timestamp 1711653199
transform 1 0 2900 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5416
timestamp 1711653199
transform 1 0 2484 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_5417
timestamp 1711653199
transform 1 0 2940 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5418
timestamp 1711653199
transform 1 0 2892 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_5419
timestamp 1711653199
transform 1 0 2916 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_5420
timestamp 1711653199
transform 1 0 2852 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_5421
timestamp 1711653199
transform 1 0 2900 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5422
timestamp 1711653199
transform 1 0 2884 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_5423
timestamp 1711653199
transform 1 0 2820 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5424
timestamp 1711653199
transform 1 0 2820 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5425
timestamp 1711653199
transform 1 0 2940 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5426
timestamp 1711653199
transform 1 0 2724 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5427
timestamp 1711653199
transform 1 0 2788 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5428
timestamp 1711653199
transform 1 0 2772 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5429
timestamp 1711653199
transform 1 0 2756 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5430
timestamp 1711653199
transform 1 0 2452 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5431
timestamp 1711653199
transform 1 0 2516 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5432
timestamp 1711653199
transform 1 0 2484 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5433
timestamp 1711653199
transform 1 0 2940 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5434
timestamp 1711653199
transform 1 0 2860 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5435
timestamp 1711653199
transform 1 0 2868 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5436
timestamp 1711653199
transform 1 0 2764 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5437
timestamp 1711653199
transform 1 0 2404 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5438
timestamp 1711653199
transform 1 0 2940 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5439
timestamp 1711653199
transform 1 0 2740 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5440
timestamp 1711653199
transform 1 0 2700 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5441
timestamp 1711653199
transform 1 0 2420 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5442
timestamp 1711653199
transform 1 0 3316 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5443
timestamp 1711653199
transform 1 0 3140 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5444
timestamp 1711653199
transform 1 0 3132 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5445
timestamp 1711653199
transform 1 0 3132 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5446
timestamp 1711653199
transform 1 0 3084 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5447
timestamp 1711653199
transform 1 0 3036 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5448
timestamp 1711653199
transform 1 0 2996 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5449
timestamp 1711653199
transform 1 0 3116 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5450
timestamp 1711653199
transform 1 0 2940 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_5451
timestamp 1711653199
transform 1 0 2916 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_5452
timestamp 1711653199
transform 1 0 2444 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_5453
timestamp 1711653199
transform 1 0 3108 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5454
timestamp 1711653199
transform 1 0 3076 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5455
timestamp 1711653199
transform 1 0 3076 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5456
timestamp 1711653199
transform 1 0 3036 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5457
timestamp 1711653199
transform 1 0 3084 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5458
timestamp 1711653199
transform 1 0 3020 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_5459
timestamp 1711653199
transform 1 0 3068 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_5460
timestamp 1711653199
transform 1 0 2948 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_5461
timestamp 1711653199
transform 1 0 3132 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5462
timestamp 1711653199
transform 1 0 3132 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5463
timestamp 1711653199
transform 1 0 3092 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5464
timestamp 1711653199
transform 1 0 3084 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5465
timestamp 1711653199
transform 1 0 3052 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5466
timestamp 1711653199
transform 1 0 3020 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5467
timestamp 1711653199
transform 1 0 3060 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5468
timestamp 1711653199
transform 1 0 2940 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5469
timestamp 1711653199
transform 1 0 3100 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5470
timestamp 1711653199
transform 1 0 2972 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5471
timestamp 1711653199
transform 1 0 3052 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5472
timestamp 1711653199
transform 1 0 2956 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5473
timestamp 1711653199
transform 1 0 3012 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5474
timestamp 1711653199
transform 1 0 2956 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5475
timestamp 1711653199
transform 1 0 2820 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5476
timestamp 1711653199
transform 1 0 3092 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5477
timestamp 1711653199
transform 1 0 3020 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_5478
timestamp 1711653199
transform 1 0 3020 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_5479
timestamp 1711653199
transform 1 0 2988 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_5480
timestamp 1711653199
transform 1 0 3356 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5481
timestamp 1711653199
transform 1 0 3324 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_5482
timestamp 1711653199
transform 1 0 3332 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_5483
timestamp 1711653199
transform 1 0 3292 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5484
timestamp 1711653199
transform 1 0 3292 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_5485
timestamp 1711653199
transform 1 0 3188 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5486
timestamp 1711653199
transform 1 0 3364 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5487
timestamp 1711653199
transform 1 0 3356 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5488
timestamp 1711653199
transform 1 0 3332 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5489
timestamp 1711653199
transform 1 0 3332 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5490
timestamp 1711653199
transform 1 0 3348 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_5491
timestamp 1711653199
transform 1 0 3348 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_5492
timestamp 1711653199
transform 1 0 3308 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5493
timestamp 1711653199
transform 1 0 3308 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_5494
timestamp 1711653199
transform 1 0 3308 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_5495
timestamp 1711653199
transform 1 0 3276 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5496
timestamp 1711653199
transform 1 0 3380 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5497
timestamp 1711653199
transform 1 0 3364 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5498
timestamp 1711653199
transform 1 0 3388 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5499
timestamp 1711653199
transform 1 0 3332 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5500
timestamp 1711653199
transform 1 0 3252 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5501
timestamp 1711653199
transform 1 0 3156 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5502
timestamp 1711653199
transform 1 0 3076 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5503
timestamp 1711653199
transform 1 0 2892 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5504
timestamp 1711653199
transform 1 0 2748 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5505
timestamp 1711653199
transform 1 0 3284 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5506
timestamp 1711653199
transform 1 0 3172 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5507
timestamp 1711653199
transform 1 0 3108 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5508
timestamp 1711653199
transform 1 0 2908 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5509
timestamp 1711653199
transform 1 0 2780 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5510
timestamp 1711653199
transform 1 0 3332 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_5511
timestamp 1711653199
transform 1 0 3300 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_5512
timestamp 1711653199
transform 1 0 3324 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5513
timestamp 1711653199
transform 1 0 3244 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5514
timestamp 1711653199
transform 1 0 3348 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_5515
timestamp 1711653199
transform 1 0 3180 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_5516
timestamp 1711653199
transform 1 0 3260 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5517
timestamp 1711653199
transform 1 0 3180 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_5518
timestamp 1711653199
transform 1 0 3252 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_5519
timestamp 1711653199
transform 1 0 3212 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_5520
timestamp 1711653199
transform 1 0 3260 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5521
timestamp 1711653199
transform 1 0 3188 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_5522
timestamp 1711653199
transform 1 0 3268 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5523
timestamp 1711653199
transform 1 0 3188 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_5524
timestamp 1711653199
transform 1 0 2796 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5525
timestamp 1711653199
transform 1 0 2684 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_5526
timestamp 1711653199
transform 1 0 2444 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5527
timestamp 1711653199
transform 1 0 2420 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5528
timestamp 1711653199
transform 1 0 2316 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5529
timestamp 1711653199
transform 1 0 2212 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5530
timestamp 1711653199
transform 1 0 2740 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5531
timestamp 1711653199
transform 1 0 2636 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5532
timestamp 1711653199
transform 1 0 964 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5533
timestamp 1711653199
transform 1 0 868 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5534
timestamp 1711653199
transform 1 0 788 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5535
timestamp 1711653199
transform 1 0 628 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5536
timestamp 1711653199
transform 1 0 1108 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5537
timestamp 1711653199
transform 1 0 1044 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5538
timestamp 1711653199
transform 1 0 452 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5539
timestamp 1711653199
transform 1 0 404 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5540
timestamp 1711653199
transform 1 0 404 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5541
timestamp 1711653199
transform 1 0 308 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5542
timestamp 1711653199
transform 1 0 220 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5543
timestamp 1711653199
transform 1 0 140 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5544
timestamp 1711653199
transform 1 0 220 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5545
timestamp 1711653199
transform 1 0 132 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5546
timestamp 1711653199
transform 1 0 180 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5547
timestamp 1711653199
transform 1 0 132 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5548
timestamp 1711653199
transform 1 0 500 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5549
timestamp 1711653199
transform 1 0 468 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5550
timestamp 1711653199
transform 1 0 2644 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5551
timestamp 1711653199
transform 1 0 2580 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5552
timestamp 1711653199
transform 1 0 2716 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5553
timestamp 1711653199
transform 1 0 2628 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5554
timestamp 1711653199
transform 1 0 2556 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5555
timestamp 1711653199
transform 1 0 2540 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5556
timestamp 1711653199
transform 1 0 2484 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5557
timestamp 1711653199
transform 1 0 2404 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5558
timestamp 1711653199
transform 1 0 2380 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5559
timestamp 1711653199
transform 1 0 2380 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5560
timestamp 1711653199
transform 1 0 2404 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5561
timestamp 1711653199
transform 1 0 2372 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5562
timestamp 1711653199
transform 1 0 2540 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5563
timestamp 1711653199
transform 1 0 2508 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5564
timestamp 1711653199
transform 1 0 2516 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5565
timestamp 1711653199
transform 1 0 2268 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5566
timestamp 1711653199
transform 1 0 2244 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5567
timestamp 1711653199
transform 1 0 2108 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5568
timestamp 1711653199
transform 1 0 2084 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5569
timestamp 1711653199
transform 1 0 2012 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5570
timestamp 1711653199
transform 1 0 1684 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5571
timestamp 1711653199
transform 1 0 2396 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5572
timestamp 1711653199
transform 1 0 2244 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5573
timestamp 1711653199
transform 1 0 2612 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5574
timestamp 1711653199
transform 1 0 2444 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5575
timestamp 1711653199
transform 1 0 2468 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5576
timestamp 1711653199
transform 1 0 2348 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5577
timestamp 1711653199
transform 1 0 2228 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5578
timestamp 1711653199
transform 1 0 2204 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5579
timestamp 1711653199
transform 1 0 2204 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5580
timestamp 1711653199
transform 1 0 1516 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5581
timestamp 1711653199
transform 1 0 2284 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5582
timestamp 1711653199
transform 1 0 2180 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5583
timestamp 1711653199
transform 1 0 2172 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5584
timestamp 1711653199
transform 1 0 1380 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5585
timestamp 1711653199
transform 1 0 2388 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5586
timestamp 1711653199
transform 1 0 2316 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5587
timestamp 1711653199
transform 1 0 2396 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5588
timestamp 1711653199
transform 1 0 2364 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5589
timestamp 1711653199
transform 1 0 2236 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5590
timestamp 1711653199
transform 1 0 2124 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5591
timestamp 1711653199
transform 1 0 1980 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5592
timestamp 1711653199
transform 1 0 3124 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5593
timestamp 1711653199
transform 1 0 2732 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5594
timestamp 1711653199
transform 1 0 2692 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5595
timestamp 1711653199
transform 1 0 2652 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5596
timestamp 1711653199
transform 1 0 1388 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5597
timestamp 1711653199
transform 1 0 1180 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5598
timestamp 1711653199
transform 1 0 1100 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5599
timestamp 1711653199
transform 1 0 1044 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5600
timestamp 1711653199
transform 1 0 1132 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5601
timestamp 1711653199
transform 1 0 1108 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5602
timestamp 1711653199
transform 1 0 964 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5603
timestamp 1711653199
transform 1 0 916 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5604
timestamp 1711653199
transform 1 0 852 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5605
timestamp 1711653199
transform 1 0 1268 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5606
timestamp 1711653199
transform 1 0 1252 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5607
timestamp 1711653199
transform 1 0 1212 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5608
timestamp 1711653199
transform 1 0 1188 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5609
timestamp 1711653199
transform 1 0 1180 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5610
timestamp 1711653199
transform 1 0 1396 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5611
timestamp 1711653199
transform 1 0 1308 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5612
timestamp 1711653199
transform 1 0 1252 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5613
timestamp 1711653199
transform 1 0 1164 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5614
timestamp 1711653199
transform 1 0 1500 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_5615
timestamp 1711653199
transform 1 0 1404 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_5616
timestamp 1711653199
transform 1 0 1332 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_5617
timestamp 1711653199
transform 1 0 1324 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5618
timestamp 1711653199
transform 1 0 1276 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5619
timestamp 1711653199
transform 1 0 1276 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5620
timestamp 1711653199
transform 1 0 1204 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5621
timestamp 1711653199
transform 1 0 1204 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5622
timestamp 1711653199
transform 1 0 900 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5623
timestamp 1711653199
transform 1 0 780 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5624
timestamp 1711653199
transform 1 0 1660 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5625
timestamp 1711653199
transform 1 0 1524 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5626
timestamp 1711653199
transform 1 0 1364 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5627
timestamp 1711653199
transform 1 0 1884 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5628
timestamp 1711653199
transform 1 0 1796 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5629
timestamp 1711653199
transform 1 0 1732 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5630
timestamp 1711653199
transform 1 0 1668 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5631
timestamp 1711653199
transform 1 0 1588 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5632
timestamp 1711653199
transform 1 0 1540 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5633
timestamp 1711653199
transform 1 0 1460 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5634
timestamp 1711653199
transform 1 0 1332 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5635
timestamp 1711653199
transform 1 0 1780 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5636
timestamp 1711653199
transform 1 0 1644 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5637
timestamp 1711653199
transform 1 0 1836 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5638
timestamp 1711653199
transform 1 0 1708 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_5639
timestamp 1711653199
transform 1 0 1572 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5640
timestamp 1711653199
transform 1 0 1492 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5641
timestamp 1711653199
transform 1 0 1524 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5642
timestamp 1711653199
transform 1 0 1492 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_5643
timestamp 1711653199
transform 1 0 1524 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5644
timestamp 1711653199
transform 1 0 1436 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5645
timestamp 1711653199
transform 1 0 1340 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5646
timestamp 1711653199
transform 1 0 1228 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5647
timestamp 1711653199
transform 1 0 1972 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5648
timestamp 1711653199
transform 1 0 1484 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5649
timestamp 1711653199
transform 1 0 1444 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5650
timestamp 1711653199
transform 1 0 1316 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5651
timestamp 1711653199
transform 1 0 1388 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5652
timestamp 1711653199
transform 1 0 1252 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5653
timestamp 1711653199
transform 1 0 1244 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5654
timestamp 1711653199
transform 1 0 1092 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5655
timestamp 1711653199
transform 1 0 1508 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5656
timestamp 1711653199
transform 1 0 1396 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5657
timestamp 1711653199
transform 1 0 1404 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5658
timestamp 1711653199
transform 1 0 1268 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5659
timestamp 1711653199
transform 1 0 1164 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5660
timestamp 1711653199
transform 1 0 1028 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5661
timestamp 1711653199
transform 1 0 964 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5662
timestamp 1711653199
transform 1 0 1404 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5663
timestamp 1711653199
transform 1 0 1348 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5664
timestamp 1711653199
transform 1 0 1332 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5665
timestamp 1711653199
transform 1 0 1308 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5666
timestamp 1711653199
transform 1 0 1356 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5667
timestamp 1711653199
transform 1 0 1324 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5668
timestamp 1711653199
transform 1 0 1228 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5669
timestamp 1711653199
transform 1 0 1084 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5670
timestamp 1711653199
transform 1 0 996 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5671
timestamp 1711653199
transform 1 0 1252 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5672
timestamp 1711653199
transform 1 0 1076 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_5673
timestamp 1711653199
transform 1 0 1004 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5674
timestamp 1711653199
transform 1 0 956 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5675
timestamp 1711653199
transform 1 0 1236 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5676
timestamp 1711653199
transform 1 0 988 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5677
timestamp 1711653199
transform 1 0 1220 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5678
timestamp 1711653199
transform 1 0 1188 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5679
timestamp 1711653199
transform 1 0 1380 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5680
timestamp 1711653199
transform 1 0 1196 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_5681
timestamp 1711653199
transform 1 0 1180 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5682
timestamp 1711653199
transform 1 0 1156 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5683
timestamp 1711653199
transform 1 0 1156 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5684
timestamp 1711653199
transform 1 0 1108 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5685
timestamp 1711653199
transform 1 0 1012 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5686
timestamp 1711653199
transform 1 0 1036 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5687
timestamp 1711653199
transform 1 0 892 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5688
timestamp 1711653199
transform 1 0 892 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5689
timestamp 1711653199
transform 1 0 868 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5690
timestamp 1711653199
transform 1 0 1100 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5691
timestamp 1711653199
transform 1 0 828 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5692
timestamp 1711653199
transform 1 0 828 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5693
timestamp 1711653199
transform 1 0 764 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5694
timestamp 1711653199
transform 1 0 732 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5695
timestamp 1711653199
transform 1 0 692 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5696
timestamp 1711653199
transform 1 0 716 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5697
timestamp 1711653199
transform 1 0 604 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_5698
timestamp 1711653199
transform 1 0 1012 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5699
timestamp 1711653199
transform 1 0 836 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5700
timestamp 1711653199
transform 1 0 636 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5701
timestamp 1711653199
transform 1 0 628 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5702
timestamp 1711653199
transform 1 0 564 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5703
timestamp 1711653199
transform 1 0 852 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5704
timestamp 1711653199
transform 1 0 676 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5705
timestamp 1711653199
transform 1 0 796 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5706
timestamp 1711653199
transform 1 0 596 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_5707
timestamp 1711653199
transform 1 0 452 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5708
timestamp 1711653199
transform 1 0 380 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5709
timestamp 1711653199
transform 1 0 556 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5710
timestamp 1711653199
transform 1 0 476 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5711
timestamp 1711653199
transform 1 0 700 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5712
timestamp 1711653199
transform 1 0 556 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5713
timestamp 1711653199
transform 1 0 404 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5714
timestamp 1711653199
transform 1 0 300 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_5715
timestamp 1711653199
transform 1 0 588 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5716
timestamp 1711653199
transform 1 0 444 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_5717
timestamp 1711653199
transform 1 0 740 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5718
timestamp 1711653199
transform 1 0 620 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5719
timestamp 1711653199
transform 1 0 948 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5720
timestamp 1711653199
transform 1 0 868 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5721
timestamp 1711653199
transform 1 0 844 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_5722
timestamp 1711653199
transform 1 0 884 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5723
timestamp 1711653199
transform 1 0 636 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5724
timestamp 1711653199
transform 1 0 524 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5725
timestamp 1711653199
transform 1 0 980 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5726
timestamp 1711653199
transform 1 0 836 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5727
timestamp 1711653199
transform 1 0 828 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5728
timestamp 1711653199
transform 1 0 716 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5729
timestamp 1711653199
transform 1 0 668 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5730
timestamp 1711653199
transform 1 0 636 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5731
timestamp 1711653199
transform 1 0 620 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5732
timestamp 1711653199
transform 1 0 620 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5733
timestamp 1711653199
transform 1 0 236 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_5734
timestamp 1711653199
transform 1 0 676 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5735
timestamp 1711653199
transform 1 0 612 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_5736
timestamp 1711653199
transform 1 0 860 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_5737
timestamp 1711653199
transform 1 0 844 0 1 2875
box -3 -3 3 3
use M3_M2  M3_M2_5738
timestamp 1711653199
transform 1 0 844 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_5739
timestamp 1711653199
transform 1 0 756 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_5740
timestamp 1711653199
transform 1 0 692 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_5741
timestamp 1711653199
transform 1 0 564 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5742
timestamp 1711653199
transform 1 0 436 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_5743
timestamp 1711653199
transform 1 0 636 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5744
timestamp 1711653199
transform 1 0 540 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5745
timestamp 1711653199
transform 1 0 476 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_5746
timestamp 1711653199
transform 1 0 244 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_5747
timestamp 1711653199
transform 1 0 476 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5748
timestamp 1711653199
transform 1 0 428 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5749
timestamp 1711653199
transform 1 0 676 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5750
timestamp 1711653199
transform 1 0 460 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_5751
timestamp 1711653199
transform 1 0 516 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5752
timestamp 1711653199
transform 1 0 260 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5753
timestamp 1711653199
transform 1 0 740 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5754
timestamp 1711653199
transform 1 0 492 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5755
timestamp 1711653199
transform 1 0 1060 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5756
timestamp 1711653199
transform 1 0 1028 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5757
timestamp 1711653199
transform 1 0 988 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5758
timestamp 1711653199
transform 1 0 972 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5759
timestamp 1711653199
transform 1 0 948 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5760
timestamp 1711653199
transform 1 0 852 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5761
timestamp 1711653199
transform 1 0 1092 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5762
timestamp 1711653199
transform 1 0 940 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5763
timestamp 1711653199
transform 1 0 908 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5764
timestamp 1711653199
transform 1 0 1172 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5765
timestamp 1711653199
transform 1 0 988 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5766
timestamp 1711653199
transform 1 0 892 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5767
timestamp 1711653199
transform 1 0 588 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5768
timestamp 1711653199
transform 1 0 572 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5769
timestamp 1711653199
transform 1 0 692 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5770
timestamp 1711653199
transform 1 0 628 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5771
timestamp 1711653199
transform 1 0 1012 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5772
timestamp 1711653199
transform 1 0 716 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5773
timestamp 1711653199
transform 1 0 1220 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5774
timestamp 1711653199
transform 1 0 1012 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5775
timestamp 1711653199
transform 1 0 932 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_5776
timestamp 1711653199
transform 1 0 932 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5777
timestamp 1711653199
transform 1 0 836 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_5778
timestamp 1711653199
transform 1 0 836 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5779
timestamp 1711653199
transform 1 0 796 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5780
timestamp 1711653199
transform 1 0 572 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5781
timestamp 1711653199
transform 1 0 404 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5782
timestamp 1711653199
transform 1 0 668 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5783
timestamp 1711653199
transform 1 0 604 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5784
timestamp 1711653199
transform 1 0 804 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_5785
timestamp 1711653199
transform 1 0 668 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5786
timestamp 1711653199
transform 1 0 844 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5787
timestamp 1711653199
transform 1 0 748 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5788
timestamp 1711653199
transform 1 0 956 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5789
timestamp 1711653199
transform 1 0 908 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_5790
timestamp 1711653199
transform 1 0 940 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5791
timestamp 1711653199
transform 1 0 916 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_5792
timestamp 1711653199
transform 1 0 1316 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5793
timestamp 1711653199
transform 1 0 1252 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_5794
timestamp 1711653199
transform 1 0 1252 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5795
timestamp 1711653199
transform 1 0 1196 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5796
timestamp 1711653199
transform 1 0 1084 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5797
timestamp 1711653199
transform 1 0 1060 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5798
timestamp 1711653199
transform 1 0 1292 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_5799
timestamp 1711653199
transform 1 0 1220 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_5800
timestamp 1711653199
transform 1 0 1116 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_5801
timestamp 1711653199
transform 1 0 1100 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_5802
timestamp 1711653199
transform 1 0 1068 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_5803
timestamp 1711653199
transform 1 0 1228 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5804
timestamp 1711653199
transform 1 0 1140 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5805
timestamp 1711653199
transform 1 0 1420 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5806
timestamp 1711653199
transform 1 0 1060 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5807
timestamp 1711653199
transform 1 0 1692 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5808
timestamp 1711653199
transform 1 0 1604 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_5809
timestamp 1711653199
transform 1 0 1468 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_5810
timestamp 1711653199
transform 1 0 1260 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_5811
timestamp 1711653199
transform 1 0 1596 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5812
timestamp 1711653199
transform 1 0 1532 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5813
timestamp 1711653199
transform 1 0 1516 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5814
timestamp 1711653199
transform 1 0 1108 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_5815
timestamp 1711653199
transform 1 0 1764 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5816
timestamp 1711653199
transform 1 0 1684 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5817
timestamp 1711653199
transform 1 0 1660 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_5818
timestamp 1711653199
transform 1 0 1212 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_5819
timestamp 1711653199
transform 1 0 1860 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5820
timestamp 1711653199
transform 1 0 1700 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5821
timestamp 1711653199
transform 1 0 1660 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5822
timestamp 1711653199
transform 1 0 1284 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_5823
timestamp 1711653199
transform 1 0 1692 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5824
timestamp 1711653199
transform 1 0 1300 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5825
timestamp 1711653199
transform 1 0 1236 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5826
timestamp 1711653199
transform 1 0 1164 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5827
timestamp 1711653199
transform 1 0 1276 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5828
timestamp 1711653199
transform 1 0 1228 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5829
timestamp 1711653199
transform 1 0 1164 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_5830
timestamp 1711653199
transform 1 0 1468 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5831
timestamp 1711653199
transform 1 0 1284 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_5832
timestamp 1711653199
transform 1 0 1716 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5833
timestamp 1711653199
transform 1 0 1692 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5834
timestamp 1711653199
transform 1 0 2740 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5835
timestamp 1711653199
transform 1 0 2652 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5836
timestamp 1711653199
transform 1 0 2188 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5837
timestamp 1711653199
transform 1 0 2140 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_5838
timestamp 1711653199
transform 1 0 2548 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5839
timestamp 1711653199
transform 1 0 2460 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5840
timestamp 1711653199
transform 1 0 1492 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5841
timestamp 1711653199
transform 1 0 1452 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5842
timestamp 1711653199
transform 1 0 716 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5843
timestamp 1711653199
transform 1 0 628 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5844
timestamp 1711653199
transform 1 0 340 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5845
timestamp 1711653199
transform 1 0 300 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_5846
timestamp 1711653199
transform 1 0 420 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5847
timestamp 1711653199
transform 1 0 356 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_5848
timestamp 1711653199
transform 1 0 244 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5849
timestamp 1711653199
transform 1 0 140 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_5850
timestamp 1711653199
transform 1 0 244 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5851
timestamp 1711653199
transform 1 0 132 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5852
timestamp 1711653199
transform 1 0 556 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5853
timestamp 1711653199
transform 1 0 468 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5854
timestamp 1711653199
transform 1 0 396 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5855
timestamp 1711653199
transform 1 0 324 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5856
timestamp 1711653199
transform 1 0 716 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5857
timestamp 1711653199
transform 1 0 604 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5858
timestamp 1711653199
transform 1 0 932 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5859
timestamp 1711653199
transform 1 0 836 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_5860
timestamp 1711653199
transform 1 0 1412 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5861
timestamp 1711653199
transform 1 0 1316 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5862
timestamp 1711653199
transform 1 0 2988 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5863
timestamp 1711653199
transform 1 0 2852 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_5864
timestamp 1711653199
transform 1 0 3356 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5865
timestamp 1711653199
transform 1 0 3252 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_5866
timestamp 1711653199
transform 1 0 3316 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5867
timestamp 1711653199
transform 1 0 3292 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_5868
timestamp 1711653199
transform 1 0 3316 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5869
timestamp 1711653199
transform 1 0 3212 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_5870
timestamp 1711653199
transform 1 0 3244 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5871
timestamp 1711653199
transform 1 0 3212 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5872
timestamp 1711653199
transform 1 0 3076 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5873
timestamp 1711653199
transform 1 0 3052 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_5874
timestamp 1711653199
transform 1 0 3284 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5875
timestamp 1711653199
transform 1 0 3220 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_5876
timestamp 1711653199
transform 1 0 3236 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5877
timestamp 1711653199
transform 1 0 3204 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5878
timestamp 1711653199
transform 1 0 3260 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5879
timestamp 1711653199
transform 1 0 3244 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5880
timestamp 1711653199
transform 1 0 3140 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5881
timestamp 1711653199
transform 1 0 3092 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_5882
timestamp 1711653199
transform 1 0 3068 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5883
timestamp 1711653199
transform 1 0 2980 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5884
timestamp 1711653199
transform 1 0 3212 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5885
timestamp 1711653199
transform 1 0 3108 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_5886
timestamp 1711653199
transform 1 0 3196 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5887
timestamp 1711653199
transform 1 0 2996 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5888
timestamp 1711653199
transform 1 0 3284 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5889
timestamp 1711653199
transform 1 0 3228 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5890
timestamp 1711653199
transform 1 0 3100 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5891
timestamp 1711653199
transform 1 0 3028 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5892
timestamp 1711653199
transform 1 0 3028 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5893
timestamp 1711653199
transform 1 0 2852 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_5894
timestamp 1711653199
transform 1 0 2852 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_5895
timestamp 1711653199
transform 1 0 2828 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5896
timestamp 1711653199
transform 1 0 2796 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_5897
timestamp 1711653199
transform 1 0 1596 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5898
timestamp 1711653199
transform 1 0 1380 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5899
timestamp 1711653199
transform 1 0 1372 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5900
timestamp 1711653199
transform 1 0 1340 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5901
timestamp 1711653199
transform 1 0 1076 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_5902
timestamp 1711653199
transform 1 0 3060 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5903
timestamp 1711653199
transform 1 0 2676 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5904
timestamp 1711653199
transform 1 0 2572 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5905
timestamp 1711653199
transform 1 0 2388 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5906
timestamp 1711653199
transform 1 0 2340 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_5907
timestamp 1711653199
transform 1 0 1924 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5908
timestamp 1711653199
transform 1 0 1924 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_5909
timestamp 1711653199
transform 1 0 1908 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_5910
timestamp 1711653199
transform 1 0 1884 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5911
timestamp 1711653199
transform 1 0 1596 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5912
timestamp 1711653199
transform 1 0 564 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_5913
timestamp 1711653199
transform 1 0 556 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_5914
timestamp 1711653199
transform 1 0 492 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5915
timestamp 1711653199
transform 1 0 428 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5916
timestamp 1711653199
transform 1 0 188 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5917
timestamp 1711653199
transform 1 0 2316 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_5918
timestamp 1711653199
transform 1 0 2316 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5919
timestamp 1711653199
transform 1 0 2268 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5920
timestamp 1711653199
transform 1 0 2228 0 1 2275
box -3 -3 3 3
use M3_M2  M3_M2_5921
timestamp 1711653199
transform 1 0 2212 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5922
timestamp 1711653199
transform 1 0 1876 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5923
timestamp 1711653199
transform 1 0 1876 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_5924
timestamp 1711653199
transform 1 0 1772 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5925
timestamp 1711653199
transform 1 0 1772 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_5926
timestamp 1711653199
transform 1 0 1756 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5927
timestamp 1711653199
transform 1 0 1300 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_5928
timestamp 1711653199
transform 1 0 1300 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5929
timestamp 1711653199
transform 1 0 1236 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_5930
timestamp 1711653199
transform 1 0 2532 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_5931
timestamp 1711653199
transform 1 0 2284 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5932
timestamp 1711653199
transform 1 0 2284 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_5933
timestamp 1711653199
transform 1 0 1924 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_5934
timestamp 1711653199
transform 1 0 1892 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5935
timestamp 1711653199
transform 1 0 1596 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5936
timestamp 1711653199
transform 1 0 1596 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_5937
timestamp 1711653199
transform 1 0 1556 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5938
timestamp 1711653199
transform 1 0 1412 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_5939
timestamp 1711653199
transform 1 0 2948 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_5940
timestamp 1711653199
transform 1 0 2828 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_5941
timestamp 1711653199
transform 1 0 2828 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_5942
timestamp 1711653199
transform 1 0 2596 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_5943
timestamp 1711653199
transform 1 0 2588 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5944
timestamp 1711653199
transform 1 0 2164 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5945
timestamp 1711653199
transform 1 0 1804 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5946
timestamp 1711653199
transform 1 0 1276 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_5947
timestamp 1711653199
transform 1 0 2844 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5948
timestamp 1711653199
transform 1 0 2844 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5949
timestamp 1711653199
transform 1 0 2828 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5950
timestamp 1711653199
transform 1 0 2692 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5951
timestamp 1711653199
transform 1 0 2684 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_5952
timestamp 1711653199
transform 1 0 2668 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_5953
timestamp 1711653199
transform 1 0 2660 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_5954
timestamp 1711653199
transform 1 0 1956 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5955
timestamp 1711653199
transform 1 0 1764 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5956
timestamp 1711653199
transform 1 0 1292 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_5957
timestamp 1711653199
transform 1 0 2596 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5958
timestamp 1711653199
transform 1 0 2580 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_5959
timestamp 1711653199
transform 1 0 2572 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_5960
timestamp 1711653199
transform 1 0 2412 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5961
timestamp 1711653199
transform 1 0 2412 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_5962
timestamp 1711653199
transform 1 0 2332 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_5963
timestamp 1711653199
transform 1 0 2308 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5964
timestamp 1711653199
transform 1 0 2132 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5965
timestamp 1711653199
transform 1 0 2132 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_5966
timestamp 1711653199
transform 1 0 1948 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5967
timestamp 1711653199
transform 1 0 1948 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_5968
timestamp 1711653199
transform 1 0 1868 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5969
timestamp 1711653199
transform 1 0 1468 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_5970
timestamp 1711653199
transform 1 0 2660 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5971
timestamp 1711653199
transform 1 0 2412 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5972
timestamp 1711653199
transform 1 0 2404 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5973
timestamp 1711653199
transform 1 0 2372 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5974
timestamp 1711653199
transform 1 0 2364 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_5975
timestamp 1711653199
transform 1 0 2324 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5976
timestamp 1711653199
transform 1 0 2324 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_5977
timestamp 1711653199
transform 1 0 2292 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_5978
timestamp 1711653199
transform 1 0 2292 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5979
timestamp 1711653199
transform 1 0 2132 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5980
timestamp 1711653199
transform 1 0 2060 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_5981
timestamp 1711653199
transform 1 0 2052 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5982
timestamp 1711653199
transform 1 0 1996 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5983
timestamp 1711653199
transform 1 0 1996 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_5984
timestamp 1711653199
transform 1 0 1572 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_5985
timestamp 1711653199
transform 1 0 2164 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_5986
timestamp 1711653199
transform 1 0 2164 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5987
timestamp 1711653199
transform 1 0 2132 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_5988
timestamp 1711653199
transform 1 0 2124 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5989
timestamp 1711653199
transform 1 0 1652 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_5990
timestamp 1711653199
transform 1 0 1636 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_5991
timestamp 1711653199
transform 1 0 2092 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5992
timestamp 1711653199
transform 1 0 2060 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5993
timestamp 1711653199
transform 1 0 2060 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5994
timestamp 1711653199
transform 1 0 2060 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5995
timestamp 1711653199
transform 1 0 2020 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5996
timestamp 1711653199
transform 1 0 2020 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5997
timestamp 1711653199
transform 1 0 1756 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_5998
timestamp 1711653199
transform 1 0 1748 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_5999
timestamp 1711653199
transform 1 0 1700 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_6000
timestamp 1711653199
transform 1 0 2564 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_6001
timestamp 1711653199
transform 1 0 2492 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_6002
timestamp 1711653199
transform 1 0 2372 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_6003
timestamp 1711653199
transform 1 0 2364 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_6004
timestamp 1711653199
transform 1 0 2268 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6005
timestamp 1711653199
transform 1 0 2268 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6006
timestamp 1711653199
transform 1 0 2196 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6007
timestamp 1711653199
transform 1 0 2172 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_6008
timestamp 1711653199
transform 1 0 2068 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6009
timestamp 1711653199
transform 1 0 1852 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_6010
timestamp 1711653199
transform 1 0 2012 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_6011
timestamp 1711653199
transform 1 0 1988 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_6012
timestamp 1711653199
transform 1 0 1972 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6013
timestamp 1711653199
transform 1 0 1940 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_6014
timestamp 1711653199
transform 1 0 1932 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_6015
timestamp 1711653199
transform 1 0 1900 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6016
timestamp 1711653199
transform 1 0 1740 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_6017
timestamp 1711653199
transform 1 0 1740 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6018
timestamp 1711653199
transform 1 0 1652 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_6019
timestamp 1711653199
transform 1 0 1876 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_6020
timestamp 1711653199
transform 1 0 1732 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_6021
timestamp 1711653199
transform 1 0 1716 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_6022
timestamp 1711653199
transform 1 0 1612 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_6023
timestamp 1711653199
transform 1 0 1492 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_6024
timestamp 1711653199
transform 1 0 1644 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_6025
timestamp 1711653199
transform 1 0 1628 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_6026
timestamp 1711653199
transform 1 0 1300 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_6027
timestamp 1711653199
transform 1 0 1444 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6028
timestamp 1711653199
transform 1 0 1364 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_6029
timestamp 1711653199
transform 1 0 1364 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_6030
timestamp 1711653199
transform 1 0 1292 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6031
timestamp 1711653199
transform 1 0 1292 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_6032
timestamp 1711653199
transform 1 0 1292 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_6033
timestamp 1711653199
transform 1 0 1204 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_6034
timestamp 1711653199
transform 1 0 1284 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_6035
timestamp 1711653199
transform 1 0 1172 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_6036
timestamp 1711653199
transform 1 0 1124 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_6037
timestamp 1711653199
transform 1 0 996 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_6038
timestamp 1711653199
transform 1 0 1132 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_6039
timestamp 1711653199
transform 1 0 1100 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_6040
timestamp 1711653199
transform 1 0 1076 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_6041
timestamp 1711653199
transform 1 0 1012 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_6042
timestamp 1711653199
transform 1 0 1268 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_6043
timestamp 1711653199
transform 1 0 1132 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_6044
timestamp 1711653199
transform 1 0 1092 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_6045
timestamp 1711653199
transform 1 0 1092 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_6046
timestamp 1711653199
transform 1 0 1012 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_6047
timestamp 1711653199
transform 1 0 1012 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_6048
timestamp 1711653199
transform 1 0 996 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_6049
timestamp 1711653199
transform 1 0 876 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_6050
timestamp 1711653199
transform 1 0 868 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_6051
timestamp 1711653199
transform 1 0 756 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_6052
timestamp 1711653199
transform 1 0 356 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_6053
timestamp 1711653199
transform 1 0 1204 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_6054
timestamp 1711653199
transform 1 0 1148 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_6055
timestamp 1711653199
transform 1 0 1148 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_6056
timestamp 1711653199
transform 1 0 732 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_6057
timestamp 1711653199
transform 1 0 564 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_6058
timestamp 1711653199
transform 1 0 564 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_6059
timestamp 1711653199
transform 1 0 516 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_6060
timestamp 1711653199
transform 1 0 404 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_6061
timestamp 1711653199
transform 1 0 404 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_6062
timestamp 1711653199
transform 1 0 260 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_6063
timestamp 1711653199
transform 1 0 244 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_6064
timestamp 1711653199
transform 1 0 1076 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_6065
timestamp 1711653199
transform 1 0 636 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_6066
timestamp 1711653199
transform 1 0 636 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_6067
timestamp 1711653199
transform 1 0 268 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_6068
timestamp 1711653199
transform 1 0 228 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_6069
timestamp 1711653199
transform 1 0 1044 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_6070
timestamp 1711653199
transform 1 0 708 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_6071
timestamp 1711653199
transform 1 0 676 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_6072
timestamp 1711653199
transform 1 0 388 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_6073
timestamp 1711653199
transform 1 0 132 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_6074
timestamp 1711653199
transform 1 0 100 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_6075
timestamp 1711653199
transform 1 0 2676 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_6076
timestamp 1711653199
transform 1 0 2676 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_6077
timestamp 1711653199
transform 1 0 2628 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_6078
timestamp 1711653199
transform 1 0 2628 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_6079
timestamp 1711653199
transform 1 0 2452 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_6080
timestamp 1711653199
transform 1 0 2452 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_6081
timestamp 1711653199
transform 1 0 2388 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6082
timestamp 1711653199
transform 1 0 2380 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_6083
timestamp 1711653199
transform 1 0 2372 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_6084
timestamp 1711653199
transform 1 0 2340 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_6085
timestamp 1711653199
transform 1 0 2332 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6086
timestamp 1711653199
transform 1 0 2140 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_6087
timestamp 1711653199
transform 1 0 1796 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_6088
timestamp 1711653199
transform 1 0 748 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6089
timestamp 1711653199
transform 1 0 604 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_6090
timestamp 1711653199
transform 1 0 572 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6091
timestamp 1711653199
transform 1 0 532 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_6092
timestamp 1711653199
transform 1 0 524 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6093
timestamp 1711653199
transform 1 0 492 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_6094
timestamp 1711653199
transform 1 0 484 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_6095
timestamp 1711653199
transform 1 0 484 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6096
timestamp 1711653199
transform 1 0 700 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_6097
timestamp 1711653199
transform 1 0 604 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_6098
timestamp 1711653199
transform 1 0 516 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_6099
timestamp 1711653199
transform 1 0 492 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_6100
timestamp 1711653199
transform 1 0 492 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_6101
timestamp 1711653199
transform 1 0 484 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_6102
timestamp 1711653199
transform 1 0 444 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_6103
timestamp 1711653199
transform 1 0 444 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_6104
timestamp 1711653199
transform 1 0 428 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_6105
timestamp 1711653199
transform 1 0 420 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_6106
timestamp 1711653199
transform 1 0 788 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_6107
timestamp 1711653199
transform 1 0 756 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_6108
timestamp 1711653199
transform 1 0 580 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6109
timestamp 1711653199
transform 1 0 580 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_6110
timestamp 1711653199
transform 1 0 556 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6111
timestamp 1711653199
transform 1 0 556 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_6112
timestamp 1711653199
transform 1 0 548 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_6113
timestamp 1711653199
transform 1 0 540 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_6114
timestamp 1711653199
transform 1 0 1004 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_6115
timestamp 1711653199
transform 1 0 988 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_6116
timestamp 1711653199
transform 1 0 948 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_6117
timestamp 1711653199
transform 1 0 876 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6118
timestamp 1711653199
transform 1 0 876 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_6119
timestamp 1711653199
transform 1 0 772 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6120
timestamp 1711653199
transform 1 0 652 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_6121
timestamp 1711653199
transform 1 0 1212 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_6122
timestamp 1711653199
transform 1 0 940 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_6123
timestamp 1711653199
transform 1 0 916 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_6124
timestamp 1711653199
transform 1 0 812 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_6125
timestamp 1711653199
transform 1 0 804 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_6126
timestamp 1711653199
transform 1 0 772 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6127
timestamp 1711653199
transform 1 0 716 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6128
timestamp 1711653199
transform 1 0 716 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_6129
timestamp 1711653199
transform 1 0 988 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6130
timestamp 1711653199
transform 1 0 724 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_6131
timestamp 1711653199
transform 1 0 660 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6132
timestamp 1711653199
transform 1 0 660 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_6133
timestamp 1711653199
transform 1 0 660 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6134
timestamp 1711653199
transform 1 0 636 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_6135
timestamp 1711653199
transform 1 0 620 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_6136
timestamp 1711653199
transform 1 0 604 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6137
timestamp 1711653199
transform 1 0 1076 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_6138
timestamp 1711653199
transform 1 0 812 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_6139
timestamp 1711653199
transform 1 0 812 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_6140
timestamp 1711653199
transform 1 0 724 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_6141
timestamp 1711653199
transform 1 0 612 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_6142
timestamp 1711653199
transform 1 0 1468 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_6143
timestamp 1711653199
transform 1 0 1428 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_6144
timestamp 1711653199
transform 1 0 1348 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6145
timestamp 1711653199
transform 1 0 1340 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_6146
timestamp 1711653199
transform 1 0 1316 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6147
timestamp 1711653199
transform 1 0 932 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_6148
timestamp 1711653199
transform 1 0 924 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_6149
timestamp 1711653199
transform 1 0 924 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_6150
timestamp 1711653199
transform 1 0 876 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_6151
timestamp 1711653199
transform 1 0 708 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_6152
timestamp 1711653199
transform 1 0 700 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_6153
timestamp 1711653199
transform 1 0 668 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_6154
timestamp 1711653199
transform 1 0 1508 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6155
timestamp 1711653199
transform 1 0 1500 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_6156
timestamp 1711653199
transform 1 0 1420 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6157
timestamp 1711653199
transform 1 0 1332 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_6158
timestamp 1711653199
transform 1 0 1164 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6159
timestamp 1711653199
transform 1 0 940 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_6160
timestamp 1711653199
transform 1 0 1676 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_6161
timestamp 1711653199
transform 1 0 1644 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_6162
timestamp 1711653199
transform 1 0 1612 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_6163
timestamp 1711653199
transform 1 0 1420 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_6164
timestamp 1711653199
transform 1 0 1148 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_6165
timestamp 1711653199
transform 1 0 1148 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_6166
timestamp 1711653199
transform 1 0 964 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_6167
timestamp 1711653199
transform 1 0 2772 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_6168
timestamp 1711653199
transform 1 0 2756 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_6169
timestamp 1711653199
transform 1 0 2748 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_6170
timestamp 1711653199
transform 1 0 2420 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_6171
timestamp 1711653199
transform 1 0 2412 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_6172
timestamp 1711653199
transform 1 0 2068 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_6173
timestamp 1711653199
transform 1 0 2020 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_6174
timestamp 1711653199
transform 1 0 1980 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_6175
timestamp 1711653199
transform 1 0 1892 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6176
timestamp 1711653199
transform 1 0 3220 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6177
timestamp 1711653199
transform 1 0 3148 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6178
timestamp 1711653199
transform 1 0 2884 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6179
timestamp 1711653199
transform 1 0 3124 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6180
timestamp 1711653199
transform 1 0 2556 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6181
timestamp 1711653199
transform 1 0 2556 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_6182
timestamp 1711653199
transform 1 0 1796 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_6183
timestamp 1711653199
transform 1 0 2180 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6184
timestamp 1711653199
transform 1 0 2060 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6185
timestamp 1711653199
transform 1 0 2028 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6186
timestamp 1711653199
transform 1 0 2684 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6187
timestamp 1711653199
transform 1 0 2628 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6188
timestamp 1711653199
transform 1 0 2484 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_6189
timestamp 1711653199
transform 1 0 2628 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_6190
timestamp 1711653199
transform 1 0 2356 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6191
timestamp 1711653199
transform 1 0 2356 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_6192
timestamp 1711653199
transform 1 0 2164 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6193
timestamp 1711653199
transform 1 0 1964 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_6194
timestamp 1711653199
transform 1 0 2052 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_6195
timestamp 1711653199
transform 1 0 1964 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_6196
timestamp 1711653199
transform 1 0 1236 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_6197
timestamp 1711653199
transform 1 0 1124 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_6198
timestamp 1711653199
transform 1 0 844 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_6199
timestamp 1711653199
transform 1 0 1092 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6200
timestamp 1711653199
transform 1 0 780 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_6201
timestamp 1711653199
transform 1 0 900 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6202
timestamp 1711653199
transform 1 0 684 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_6203
timestamp 1711653199
transform 1 0 948 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6204
timestamp 1711653199
transform 1 0 724 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_6205
timestamp 1711653199
transform 1 0 820 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_6206
timestamp 1711653199
transform 1 0 780 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_6207
timestamp 1711653199
transform 1 0 860 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_6208
timestamp 1711653199
transform 1 0 820 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_6209
timestamp 1711653199
transform 1 0 756 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_6210
timestamp 1711653199
transform 1 0 956 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_6211
timestamp 1711653199
transform 1 0 804 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_6212
timestamp 1711653199
transform 1 0 764 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_6213
timestamp 1711653199
transform 1 0 1140 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_6214
timestamp 1711653199
transform 1 0 1108 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_6215
timestamp 1711653199
transform 1 0 972 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_6216
timestamp 1711653199
transform 1 0 780 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_6217
timestamp 1711653199
transform 1 0 1196 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_6218
timestamp 1711653199
transform 1 0 828 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_6219
timestamp 1711653199
transform 1 0 1308 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_6220
timestamp 1711653199
transform 1 0 1164 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_6221
timestamp 1711653199
transform 1 0 924 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_6222
timestamp 1711653199
transform 1 0 2476 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6223
timestamp 1711653199
transform 1 0 2412 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6224
timestamp 1711653199
transform 1 0 2284 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6225
timestamp 1711653199
transform 1 0 2124 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6226
timestamp 1711653199
transform 1 0 1932 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6227
timestamp 1711653199
transform 1 0 1852 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6228
timestamp 1711653199
transform 1 0 1732 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6229
timestamp 1711653199
transform 1 0 1620 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6230
timestamp 1711653199
transform 1 0 1500 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6231
timestamp 1711653199
transform 1 0 1268 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_6232
timestamp 1711653199
transform 1 0 1108 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_6233
timestamp 1711653199
transform 1 0 956 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_6234
timestamp 1711653199
transform 1 0 780 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_6235
timestamp 1711653199
transform 1 0 2716 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6236
timestamp 1711653199
transform 1 0 2692 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_6237
timestamp 1711653199
transform 1 0 2532 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6238
timestamp 1711653199
transform 1 0 2524 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_6239
timestamp 1711653199
transform 1 0 2492 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6240
timestamp 1711653199
transform 1 0 2340 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_6241
timestamp 1711653199
transform 1 0 2340 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_6242
timestamp 1711653199
transform 1 0 2220 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_6243
timestamp 1711653199
transform 1 0 2092 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_6244
timestamp 1711653199
transform 1 0 1996 0 1 3195
box -3 -3 3 3
use NAND2X1  NAND2X1_0
timestamp 1711653199
transform 1 0 2968 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_1
timestamp 1711653199
transform 1 0 2280 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_2
timestamp 1711653199
transform 1 0 1160 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_3
timestamp 1711653199
transform 1 0 288 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_4
timestamp 1711653199
transform 1 0 360 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_5
timestamp 1711653199
transform 1 0 920 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_6
timestamp 1711653199
transform 1 0 2744 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_7
timestamp 1711653199
transform 1 0 1840 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_8
timestamp 1711653199
transform 1 0 400 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_9
timestamp 1711653199
transform 1 0 2032 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_10
timestamp 1711653199
transform 1 0 1432 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_11
timestamp 1711653199
transform 1 0 1432 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_12
timestamp 1711653199
transform 1 0 1656 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_13
timestamp 1711653199
transform 1 0 384 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_14
timestamp 1711653199
transform 1 0 952 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_15
timestamp 1711653199
transform 1 0 2840 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_16
timestamp 1711653199
transform 1 0 1688 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_17
timestamp 1711653199
transform 1 0 680 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_18
timestamp 1711653199
transform 1 0 1496 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_19
timestamp 1711653199
transform 1 0 1424 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_20
timestamp 1711653199
transform 1 0 1992 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_21
timestamp 1711653199
transform 1 0 2176 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_22
timestamp 1711653199
transform 1 0 2208 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_23
timestamp 1711653199
transform 1 0 2104 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_24
timestamp 1711653199
transform 1 0 1936 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1711653199
transform 1 0 1928 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1711653199
transform 1 0 2280 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_27
timestamp 1711653199
transform 1 0 2184 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_28
timestamp 1711653199
transform 1 0 1904 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_29
timestamp 1711653199
transform 1 0 2048 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_30
timestamp 1711653199
transform 1 0 2136 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_31
timestamp 1711653199
transform 1 0 1728 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_32
timestamp 1711653199
transform 1 0 1944 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_33
timestamp 1711653199
transform 1 0 1624 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_34
timestamp 1711653199
transform 1 0 1712 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_35
timestamp 1711653199
transform 1 0 1728 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_36
timestamp 1711653199
transform 1 0 1656 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_37
timestamp 1711653199
transform 1 0 1632 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_38
timestamp 1711653199
transform 1 0 1816 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1711653199
transform 1 0 1552 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_40
timestamp 1711653199
transform 1 0 1592 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_41
timestamp 1711653199
transform 1 0 1688 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_42
timestamp 1711653199
transform 1 0 1688 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_43
timestamp 1711653199
transform 1 0 2056 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_44
timestamp 1711653199
transform 1 0 1912 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_45
timestamp 1711653199
transform 1 0 1672 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_46
timestamp 1711653199
transform 1 0 624 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_47
timestamp 1711653199
transform 1 0 768 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_48
timestamp 1711653199
transform 1 0 680 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_49
timestamp 1711653199
transform 1 0 632 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_50
timestamp 1711653199
transform 1 0 536 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_51
timestamp 1711653199
transform 1 0 752 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_52
timestamp 1711653199
transform 1 0 872 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_53
timestamp 1711653199
transform 1 0 128 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_54
timestamp 1711653199
transform 1 0 232 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_55
timestamp 1711653199
transform 1 0 248 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_56
timestamp 1711653199
transform 1 0 184 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_57
timestamp 1711653199
transform 1 0 136 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_58
timestamp 1711653199
transform 1 0 2336 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_59
timestamp 1711653199
transform 1 0 200 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_60
timestamp 1711653199
transform 1 0 336 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_61
timestamp 1711653199
transform 1 0 112 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_62
timestamp 1711653199
transform 1 0 88 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_63
timestamp 1711653199
transform 1 0 112 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_64
timestamp 1711653199
transform 1 0 136 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_65
timestamp 1711653199
transform 1 0 88 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_66
timestamp 1711653199
transform 1 0 136 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_67
timestamp 1711653199
transform 1 0 192 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_68
timestamp 1711653199
transform 1 0 2216 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_69
timestamp 1711653199
transform 1 0 88 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_70
timestamp 1711653199
transform 1 0 112 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_71
timestamp 1711653199
transform 1 0 88 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_72
timestamp 1711653199
transform 1 0 352 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_73
timestamp 1711653199
transform 1 0 400 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_74
timestamp 1711653199
transform 1 0 392 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_75
timestamp 1711653199
transform 1 0 472 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_76
timestamp 1711653199
transform 1 0 504 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_77
timestamp 1711653199
transform 1 0 128 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_78
timestamp 1711653199
transform 1 0 288 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_79
timestamp 1711653199
transform 1 0 224 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_80
timestamp 1711653199
transform 1 0 328 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_81
timestamp 1711653199
transform 1 0 312 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_82
timestamp 1711653199
transform 1 0 576 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_83
timestamp 1711653199
transform 1 0 384 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_84
timestamp 1711653199
transform 1 0 872 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_85
timestamp 1711653199
transform 1 0 384 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_86
timestamp 1711653199
transform 1 0 464 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_87
timestamp 1711653199
transform 1 0 568 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_88
timestamp 1711653199
transform 1 0 888 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_89
timestamp 1711653199
transform 1 0 696 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_90
timestamp 1711653199
transform 1 0 520 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_91
timestamp 1711653199
transform 1 0 816 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_92
timestamp 1711653199
transform 1 0 512 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_93
timestamp 1711653199
transform 1 0 1008 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_94
timestamp 1711653199
transform 1 0 1784 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_95
timestamp 1711653199
transform 1 0 2208 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_96
timestamp 1711653199
transform 1 0 1760 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_97
timestamp 1711653199
transform 1 0 1744 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_98
timestamp 1711653199
transform 1 0 976 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_99
timestamp 1711653199
transform 1 0 1832 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_100
timestamp 1711653199
transform 1 0 1672 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_101
timestamp 1711653199
transform 1 0 824 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_102
timestamp 1711653199
transform 1 0 736 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_103
timestamp 1711653199
transform 1 0 792 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_104
timestamp 1711653199
transform 1 0 944 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_105
timestamp 1711653199
transform 1 0 2592 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_106
timestamp 1711653199
transform 1 0 2328 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_107
timestamp 1711653199
transform 1 0 848 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_108
timestamp 1711653199
transform 1 0 408 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_109
timestamp 1711653199
transform 1 0 456 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_110
timestamp 1711653199
transform 1 0 432 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_111
timestamp 1711653199
transform 1 0 400 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_112
timestamp 1711653199
transform 1 0 408 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_113
timestamp 1711653199
transform 1 0 360 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_114
timestamp 1711653199
transform 1 0 512 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_115
timestamp 1711653199
transform 1 0 224 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_116
timestamp 1711653199
transform 1 0 312 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_117
timestamp 1711653199
transform 1 0 112 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_118
timestamp 1711653199
transform 1 0 192 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_119
timestamp 1711653199
transform 1 0 304 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_120
timestamp 1711653199
transform 1 0 136 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_121
timestamp 1711653199
transform 1 0 320 0 1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_122
timestamp 1711653199
transform 1 0 1368 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_123
timestamp 1711653199
transform 1 0 1248 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_124
timestamp 1711653199
transform 1 0 1280 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_125
timestamp 1711653199
transform 1 0 1392 0 -1 1970
box -8 -3 32 105
use NAND2X1  NAND2X1_126
timestamp 1711653199
transform 1 0 1432 0 -1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_127
timestamp 1711653199
transform 1 0 1296 0 1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_128
timestamp 1711653199
transform 1 0 1392 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_129
timestamp 1711653199
transform 1 0 1312 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_130
timestamp 1711653199
transform 1 0 320 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_131
timestamp 1711653199
transform 1 0 1424 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_132
timestamp 1711653199
transform 1 0 1088 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_133
timestamp 1711653199
transform 1 0 1344 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_134
timestamp 1711653199
transform 1 0 1352 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_135
timestamp 1711653199
transform 1 0 2480 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_136
timestamp 1711653199
transform 1 0 1304 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_137
timestamp 1711653199
transform 1 0 1304 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_138
timestamp 1711653199
transform 1 0 1208 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_139
timestamp 1711653199
transform 1 0 1112 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_140
timestamp 1711653199
transform 1 0 1016 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_141
timestamp 1711653199
transform 1 0 1016 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_142
timestamp 1711653199
transform 1 0 1120 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_143
timestamp 1711653199
transform 1 0 1128 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_144
timestamp 1711653199
transform 1 0 2544 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_145
timestamp 1711653199
transform 1 0 1608 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_146
timestamp 1711653199
transform 1 0 2224 0 -1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_147
timestamp 1711653199
transform 1 0 3184 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_148
timestamp 1711653199
transform 1 0 3200 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_149
timestamp 1711653199
transform 1 0 3032 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_150
timestamp 1711653199
transform 1 0 3048 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_151
timestamp 1711653199
transform 1 0 3328 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_152
timestamp 1711653199
transform 1 0 3360 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_153
timestamp 1711653199
transform 1 0 3336 0 1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_154
timestamp 1711653199
transform 1 0 3320 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_155
timestamp 1711653199
transform 1 0 3272 0 -1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_156
timestamp 1711653199
transform 1 0 3312 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_157
timestamp 1711653199
transform 1 0 3240 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_158
timestamp 1711653199
transform 1 0 3208 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_159
timestamp 1711653199
transform 1 0 3352 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_160
timestamp 1711653199
transform 1 0 3328 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_161
timestamp 1711653199
transform 1 0 3344 0 1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_162
timestamp 1711653199
transform 1 0 3248 0 1 170
box -8 -3 32 105
use NAND2X1  NAND2X1_163
timestamp 1711653199
transform 1 0 3256 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_164
timestamp 1711653199
transform 1 0 3232 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_165
timestamp 1711653199
transform 1 0 3208 0 -1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_166
timestamp 1711653199
transform 1 0 3352 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_167
timestamp 1711653199
transform 1 0 2680 0 1 370
box -8 -3 32 105
use NAND2X1  NAND2X1_168
timestamp 1711653199
transform 1 0 3000 0 -1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_169
timestamp 1711653199
transform 1 0 3168 0 1 570
box -8 -3 32 105
use NAND2X1  NAND2X1_170
timestamp 1711653199
transform 1 0 2736 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_171
timestamp 1711653199
transform 1 0 2744 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_172
timestamp 1711653199
transform 1 0 2616 0 1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_173
timestamp 1711653199
transform 1 0 2640 0 -1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_174
timestamp 1711653199
transform 1 0 3136 0 -1 1570
box -8 -3 32 105
use NAND2X1  NAND2X1_175
timestamp 1711653199
transform 1 0 2912 0 -1 2170
box -8 -3 32 105
use NAND2X1  NAND2X1_176
timestamp 1711653199
transform 1 0 2992 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_177
timestamp 1711653199
transform 1 0 2704 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_178
timestamp 1711653199
transform 1 0 3112 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_179
timestamp 1711653199
transform 1 0 3064 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_180
timestamp 1711653199
transform 1 0 3312 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_181
timestamp 1711653199
transform 1 0 3336 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_182
timestamp 1711653199
transform 1 0 3312 0 -1 2370
box -8 -3 32 105
use NAND2X1  NAND2X1_183
timestamp 1711653199
transform 1 0 3184 0 1 1770
box -8 -3 32 105
use NAND2X1  NAND2X1_184
timestamp 1711653199
transform 1 0 2656 0 1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_185
timestamp 1711653199
transform 1 0 2232 0 1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_186
timestamp 1711653199
transform 1 0 2616 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_187
timestamp 1711653199
transform 1 0 2640 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_188
timestamp 1711653199
transform 1 0 608 0 1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_189
timestamp 1711653199
transform 1 0 520 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_190
timestamp 1711653199
transform 1 0 448 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_191
timestamp 1711653199
transform 1 0 424 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_192
timestamp 1711653199
transform 1 0 600 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_193
timestamp 1711653199
transform 1 0 568 0 1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_194
timestamp 1711653199
transform 1 0 720 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_195
timestamp 1711653199
transform 1 0 936 0 -1 2570
box -8 -3 32 105
use NAND2X1  NAND2X1_196
timestamp 1711653199
transform 1 0 1248 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_197
timestamp 1711653199
transform 1 0 840 0 -1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_198
timestamp 1711653199
transform 1 0 936 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_199
timestamp 1711653199
transform 1 0 1232 0 1 2770
box -8 -3 32 105
use NAND2X1  NAND2X1_200
timestamp 1711653199
transform 1 0 3112 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_201
timestamp 1711653199
transform 1 0 3064 0 -1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_202
timestamp 1711653199
transform 1 0 3048 0 1 2770
box -8 -3 32 105
use NAND3X1  NAND3X1_0
timestamp 1711653199
transform 1 0 1536 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_1
timestamp 1711653199
transform 1 0 2384 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_2
timestamp 1711653199
transform 1 0 2392 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_3
timestamp 1711653199
transform 1 0 2520 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_4
timestamp 1711653199
transform 1 0 1736 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_5
timestamp 1711653199
transform 1 0 1152 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_6
timestamp 1711653199
transform 1 0 1608 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_7
timestamp 1711653199
transform 1 0 2368 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_8
timestamp 1711653199
transform 1 0 2592 0 -1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_9
timestamp 1711653199
transform 1 0 1640 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_10
timestamp 1711653199
transform 1 0 1536 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_11
timestamp 1711653199
transform 1 0 2752 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_12
timestamp 1711653199
transform 1 0 1800 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_13
timestamp 1711653199
transform 1 0 1992 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_14
timestamp 1711653199
transform 1 0 1896 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_15
timestamp 1711653199
transform 1 0 1592 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_16
timestamp 1711653199
transform 1 0 1888 0 -1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_17
timestamp 1711653199
transform 1 0 1816 0 1 1170
box -8 -3 40 105
use NAND3X1  NAND3X1_18
timestamp 1711653199
transform 1 0 1696 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_19
timestamp 1711653199
transform 1 0 1832 0 1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_20
timestamp 1711653199
transform 1 0 2072 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_21
timestamp 1711653199
transform 1 0 1592 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_22
timestamp 1711653199
transform 1 0 1128 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_23
timestamp 1711653199
transform 1 0 2104 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_24
timestamp 1711653199
transform 1 0 584 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_25
timestamp 1711653199
transform 1 0 592 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_26
timestamp 1711653199
transform 1 0 704 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_27
timestamp 1711653199
transform 1 0 560 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_28
timestamp 1711653199
transform 1 0 248 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_29
timestamp 1711653199
transform 1 0 224 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_30
timestamp 1711653199
transform 1 0 296 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_31
timestamp 1711653199
transform 1 0 224 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_32
timestamp 1711653199
transform 1 0 160 0 1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_33
timestamp 1711653199
transform 1 0 160 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_34
timestamp 1711653199
transform 1 0 96 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_35
timestamp 1711653199
transform 1 0 160 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_36
timestamp 1711653199
transform 1 0 448 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_37
timestamp 1711653199
transform 1 0 296 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_38
timestamp 1711653199
transform 1 0 512 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_39
timestamp 1711653199
transform 1 0 656 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_40
timestamp 1711653199
transform 1 0 488 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_41
timestamp 1711653199
transform 1 0 1008 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_42
timestamp 1711653199
transform 1 0 496 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_43
timestamp 1711653199
transform 1 0 552 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_44
timestamp 1711653199
transform 1 0 424 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_45
timestamp 1711653199
transform 1 0 640 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_46
timestamp 1711653199
transform 1 0 944 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_47
timestamp 1711653199
transform 1 0 648 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_48
timestamp 1711653199
transform 1 0 2152 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_49
timestamp 1711653199
transform 1 0 1456 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_50
timestamp 1711653199
transform 1 0 1384 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_51
timestamp 1711653199
transform 1 0 2088 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_52
timestamp 1711653199
transform 1 0 808 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_53
timestamp 1711653199
transform 1 0 736 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_54
timestamp 1711653199
transform 1 0 872 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_55
timestamp 1711653199
transform 1 0 728 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_56
timestamp 1711653199
transform 1 0 384 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_57
timestamp 1711653199
transform 1 0 392 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_58
timestamp 1711653199
transform 1 0 424 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_59
timestamp 1711653199
transform 1 0 440 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_60
timestamp 1711653199
transform 1 0 304 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_61
timestamp 1711653199
transform 1 0 248 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_62
timestamp 1711653199
transform 1 0 184 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_63
timestamp 1711653199
transform 1 0 264 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_64
timestamp 1711653199
transform 1 0 1240 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_65
timestamp 1711653199
transform 1 0 1152 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_66
timestamp 1711653199
transform 1 0 1240 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_67
timestamp 1711653199
transform 1 0 1024 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_68
timestamp 1711653199
transform 1 0 1176 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_69
timestamp 1711653199
transform 1 0 1224 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_70
timestamp 1711653199
transform 1 0 1832 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_71
timestamp 1711653199
transform 1 0 1232 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_72
timestamp 1711653199
transform 1 0 1120 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_73
timestamp 1711653199
transform 1 0 1120 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_74
timestamp 1711653199
transform 1 0 1048 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_75
timestamp 1711653199
transform 1 0 1080 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_76
timestamp 1711653199
transform 1 0 968 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_77
timestamp 1711653199
transform 1 0 2256 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_78
timestamp 1711653199
transform 1 0 2600 0 1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_79
timestamp 1711653199
transform 1 0 2520 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_80
timestamp 1711653199
transform 1 0 2304 0 1 170
box -8 -3 40 105
use NAND3X1  NAND3X1_81
timestamp 1711653199
transform 1 0 3080 0 -1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_82
timestamp 1711653199
transform 1 0 3040 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_83
timestamp 1711653199
transform 1 0 2960 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_84
timestamp 1711653199
transform 1 0 3000 0 1 1370
box -8 -3 40 105
use NAND3X1  NAND3X1_85
timestamp 1711653199
transform 1 0 3256 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_86
timestamp 1711653199
transform 1 0 3352 0 -1 570
box -8 -3 40 105
use NAND3X1  NAND3X1_87
timestamp 1711653199
transform 1 0 3344 0 1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_88
timestamp 1711653199
transform 1 0 3200 0 -1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_89
timestamp 1711653199
transform 1 0 3312 0 1 1570
box -8 -3 40 105
use NAND3X1  NAND3X1_90
timestamp 1711653199
transform 1 0 3152 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_91
timestamp 1711653199
transform 1 0 3352 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_92
timestamp 1711653199
transform 1 0 3296 0 -1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_93
timestamp 1711653199
transform 1 0 2832 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_94
timestamp 1711653199
transform 1 0 2752 0 -1 370
box -8 -3 40 105
use NAND3X1  NAND3X1_95
timestamp 1711653199
transform 1 0 1640 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_96
timestamp 1711653199
transform 1 0 2208 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_97
timestamp 1711653199
transform 1 0 2568 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_98
timestamp 1711653199
transform 1 0 2616 0 -1 1970
box -8 -3 40 105
use NAND3X1  NAND3X1_99
timestamp 1711653199
transform 1 0 2808 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_100
timestamp 1711653199
transform 1 0 2088 0 -1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_101
timestamp 1711653199
transform 1 0 2272 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_102
timestamp 1711653199
transform 1 0 2840 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_103
timestamp 1711653199
transform 1 0 2272 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_104
timestamp 1711653199
transform 1 0 2536 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_105
timestamp 1711653199
transform 1 0 2632 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_106
timestamp 1711653199
transform 1 0 2008 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_107
timestamp 1711653199
transform 1 0 2304 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_108
timestamp 1711653199
transform 1 0 2904 0 -1 970
box -8 -3 40 105
use NAND3X1  NAND3X1_109
timestamp 1711653199
transform 1 0 2976 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_110
timestamp 1711653199
transform 1 0 2352 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_111
timestamp 1711653199
transform 1 0 2736 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_112
timestamp 1711653199
transform 1 0 2904 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_113
timestamp 1711653199
transform 1 0 2424 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_114
timestamp 1711653199
transform 1 0 2912 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_115
timestamp 1711653199
transform 1 0 3000 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_116
timestamp 1711653199
transform 1 0 2856 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_117
timestamp 1711653199
transform 1 0 2384 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_118
timestamp 1711653199
transform 1 0 2224 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_119
timestamp 1711653199
transform 1 0 2872 0 -1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_120
timestamp 1711653199
transform 1 0 2192 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_121
timestamp 1711653199
transform 1 0 3352 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_122
timestamp 1711653199
transform 1 0 3320 0 -1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_123
timestamp 1711653199
transform 1 0 3208 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_124
timestamp 1711653199
transform 1 0 3240 0 -1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_125
timestamp 1711653199
transform 1 0 3352 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_126
timestamp 1711653199
transform 1 0 3312 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_127
timestamp 1711653199
transform 1 0 3304 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_128
timestamp 1711653199
transform 1 0 2656 0 1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_129
timestamp 1711653199
transform 1 0 2088 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_130
timestamp 1711653199
transform 1 0 2440 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_131
timestamp 1711653199
transform 1 0 2168 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_132
timestamp 1711653199
transform 1 0 2432 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_133
timestamp 1711653199
transform 1 0 2216 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_134
timestamp 1711653199
transform 1 0 2384 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_135
timestamp 1711653199
transform 1 0 2512 0 -1 3170
box -8 -3 40 105
use NAND3X1  NAND3X1_136
timestamp 1711653199
transform 1 0 2272 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_137
timestamp 1711653199
transform 1 0 2096 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_138
timestamp 1711653199
transform 1 0 1160 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_139
timestamp 1711653199
transform 1 0 960 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_140
timestamp 1711653199
transform 1 0 1184 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_141
timestamp 1711653199
transform 1 0 1312 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_142
timestamp 1711653199
transform 1 0 1480 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_143
timestamp 1711653199
transform 1 0 1184 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_144
timestamp 1711653199
transform 1 0 1672 0 1 2370
box -8 -3 40 105
use NAND3X1  NAND3X1_145
timestamp 1711653199
transform 1 0 1096 0 1 2570
box -8 -3 40 105
use NAND3X1  NAND3X1_146
timestamp 1711653199
transform 1 0 1112 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_147
timestamp 1711653199
transform 1 0 808 0 -1 2770
box -8 -3 40 105
use NAND3X1  NAND3X1_148
timestamp 1711653199
transform 1 0 728 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_149
timestamp 1711653199
transform 1 0 1944 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_150
timestamp 1711653199
transform 1 0 3104 0 1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_151
timestamp 1711653199
transform 1 0 3104 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_152
timestamp 1711653199
transform 1 0 3000 0 -1 2970
box -8 -3 40 105
use NAND3X1  NAND3X1_153
timestamp 1711653199
transform 1 0 3032 0 -1 2970
box -8 -3 40 105
use NOR2X1  NOR2X1_0
timestamp 1711653199
transform 1 0 2704 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_1
timestamp 1711653199
transform 1 0 2896 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_2
timestamp 1711653199
transform 1 0 2352 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_3
timestamp 1711653199
transform 1 0 2536 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_4
timestamp 1711653199
transform 1 0 1400 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1711653199
transform 1 0 1736 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_6
timestamp 1711653199
transform 1 0 1376 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_7
timestamp 1711653199
transform 1 0 1488 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_8
timestamp 1711653199
transform 1 0 2656 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_9
timestamp 1711653199
transform 1 0 1528 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_10
timestamp 1711653199
transform 1 0 1336 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_11
timestamp 1711653199
transform 1 0 1792 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_12
timestamp 1711653199
transform 1 0 1728 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_13
timestamp 1711653199
transform 1 0 1888 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_14
timestamp 1711653199
transform 1 0 528 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1711653199
transform 1 0 760 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_16
timestamp 1711653199
transform 1 0 1520 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_17
timestamp 1711653199
transform 1 0 1952 0 1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_18
timestamp 1711653199
transform 1 0 1456 0 -1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_19
timestamp 1711653199
transform 1 0 1392 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_20
timestamp 1711653199
transform 1 0 2088 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_21
timestamp 1711653199
transform 1 0 2368 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_22
timestamp 1711653199
transform 1 0 2424 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_23
timestamp 1711653199
transform 1 0 2576 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_24
timestamp 1711653199
transform 1 0 2776 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_25
timestamp 1711653199
transform 1 0 2480 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_26
timestamp 1711653199
transform 1 0 2128 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_27
timestamp 1711653199
transform 1 0 2320 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_28
timestamp 1711653199
transform 1 0 2176 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_29
timestamp 1711653199
transform 1 0 2120 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_30
timestamp 1711653199
transform 1 0 1744 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_31
timestamp 1711653199
transform 1 0 1968 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_32
timestamp 1711653199
transform 1 0 2416 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_33
timestamp 1711653199
transform 1 0 1656 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_34
timestamp 1711653199
transform 1 0 1624 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_35
timestamp 1711653199
transform 1 0 2400 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_36
timestamp 1711653199
transform 1 0 1488 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_37
timestamp 1711653199
transform 1 0 2448 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_38
timestamp 1711653199
transform 1 0 1080 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_39
timestamp 1711653199
transform 1 0 1968 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_40
timestamp 1711653199
transform 1 0 608 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_41
timestamp 1711653199
transform 1 0 2096 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_42
timestamp 1711653199
transform 1 0 2536 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_43
timestamp 1711653199
transform 1 0 2376 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_44
timestamp 1711653199
transform 1 0 712 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_45
timestamp 1711653199
transform 1 0 1552 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_46
timestamp 1711653199
transform 1 0 1520 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_47
timestamp 1711653199
transform 1 0 1608 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_48
timestamp 1711653199
transform 1 0 192 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_49
timestamp 1711653199
transform 1 0 1288 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_50
timestamp 1711653199
transform 1 0 1264 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_51
timestamp 1711653199
transform 1 0 480 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_52
timestamp 1711653199
transform 1 0 696 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_53
timestamp 1711653199
transform 1 0 864 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_54
timestamp 1711653199
transform 1 0 2240 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_55
timestamp 1711653199
transform 1 0 1224 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_56
timestamp 1711653199
transform 1 0 2080 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_57
timestamp 1711653199
transform 1 0 1648 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_58
timestamp 1711653199
transform 1 0 1480 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_59
timestamp 1711653199
transform 1 0 1496 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_60
timestamp 1711653199
transform 1 0 1440 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_61
timestamp 1711653199
transform 1 0 1968 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_62
timestamp 1711653199
transform 1 0 848 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_63
timestamp 1711653199
transform 1 0 800 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_64
timestamp 1711653199
transform 1 0 1808 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_65
timestamp 1711653199
transform 1 0 1944 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_66
timestamp 1711653199
transform 1 0 896 0 1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_67
timestamp 1711653199
transform 1 0 1560 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_68
timestamp 1711653199
transform 1 0 488 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_69
timestamp 1711653199
transform 1 0 1560 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_70
timestamp 1711653199
transform 1 0 1424 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_71
timestamp 1711653199
transform 1 0 1496 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_72
timestamp 1711653199
transform 1 0 1312 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_73
timestamp 1711653199
transform 1 0 848 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_74
timestamp 1711653199
transform 1 0 1240 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_75
timestamp 1711653199
transform 1 0 1488 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_76
timestamp 1711653199
transform 1 0 912 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_77
timestamp 1711653199
transform 1 0 864 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_78
timestamp 1711653199
transform 1 0 1176 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_79
timestamp 1711653199
transform 1 0 2104 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_80
timestamp 1711653199
transform 1 0 1616 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_81
timestamp 1711653199
transform 1 0 1880 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_82
timestamp 1711653199
transform 1 0 1728 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_83
timestamp 1711653199
transform 1 0 1072 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_84
timestamp 1711653199
transform 1 0 1656 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_85
timestamp 1711653199
transform 1 0 1536 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_86
timestamp 1711653199
transform 1 0 1232 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_87
timestamp 1711653199
transform 1 0 1472 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_88
timestamp 1711653199
transform 1 0 2272 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_89
timestamp 1711653199
transform 1 0 2392 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_90
timestamp 1711653199
transform 1 0 2040 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_91
timestamp 1711653199
transform 1 0 2152 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_92
timestamp 1711653199
transform 1 0 3160 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_93
timestamp 1711653199
transform 1 0 3184 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_94
timestamp 1711653199
transform 1 0 3112 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_95
timestamp 1711653199
transform 1 0 2920 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_96
timestamp 1711653199
transform 1 0 2248 0 -1 170
box -8 -3 32 105
use NOR2X1  NOR2X1_97
timestamp 1711653199
transform 1 0 1792 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_98
timestamp 1711653199
transform 1 0 2552 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_99
timestamp 1711653199
transform 1 0 2912 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_100
timestamp 1711653199
transform 1 0 3072 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_101
timestamp 1711653199
transform 1 0 2944 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_102
timestamp 1711653199
transform 1 0 2192 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_103
timestamp 1711653199
transform 1 0 3040 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_104
timestamp 1711653199
transform 1 0 2432 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_105
timestamp 1711653199
transform 1 0 1376 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_106
timestamp 1711653199
transform 1 0 2216 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_107
timestamp 1711653199
transform 1 0 2512 0 1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_108
timestamp 1711653199
transform 1 0 1360 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_109
timestamp 1711653199
transform 1 0 2144 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_110
timestamp 1711653199
transform 1 0 2664 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_111
timestamp 1711653199
transform 1 0 2736 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_112
timestamp 1711653199
transform 1 0 2808 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_113
timestamp 1711653199
transform 1 0 2672 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_114
timestamp 1711653199
transform 1 0 2656 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_115
timestamp 1711653199
transform 1 0 2568 0 -1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_116
timestamp 1711653199
transform 1 0 2088 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_117
timestamp 1711653199
transform 1 0 2576 0 1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_118
timestamp 1711653199
transform 1 0 2520 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_119
timestamp 1711653199
transform 1 0 2264 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_120
timestamp 1711653199
transform 1 0 2056 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_121
timestamp 1711653199
transform 1 0 2264 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_122
timestamp 1711653199
transform 1 0 2648 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_123
timestamp 1711653199
transform 1 0 2496 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_124
timestamp 1711653199
transform 1 0 2296 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_125
timestamp 1711653199
transform 1 0 2744 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_126
timestamp 1711653199
transform 1 0 2344 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_127
timestamp 1711653199
transform 1 0 2680 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_128
timestamp 1711653199
transform 1 0 2896 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_129
timestamp 1711653199
transform 1 0 2776 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_130
timestamp 1711653199
transform 1 0 2440 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_131
timestamp 1711653199
transform 1 0 2496 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_132
timestamp 1711653199
transform 1 0 2352 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_133
timestamp 1711653199
transform 1 0 2664 0 1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_134
timestamp 1711653199
transform 1 0 2800 0 -1 970
box -8 -3 32 105
use NOR2X1  NOR2X1_135
timestamp 1711653199
transform 1 0 2800 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_136
timestamp 1711653199
transform 1 0 2400 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_137
timestamp 1711653199
transform 1 0 2864 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_138
timestamp 1711653199
transform 1 0 3024 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_139
timestamp 1711653199
transform 1 0 3104 0 -1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_140
timestamp 1711653199
transform 1 0 3216 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_141
timestamp 1711653199
transform 1 0 2464 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_142
timestamp 1711653199
transform 1 0 2848 0 -1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_143
timestamp 1711653199
transform 1 0 3000 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_144
timestamp 1711653199
transform 1 0 3160 0 1 1370
box -8 -3 32 105
use NOR2X1  NOR2X1_145
timestamp 1711653199
transform 1 0 2960 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_146
timestamp 1711653199
transform 1 0 2936 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_147
timestamp 1711653199
transform 1 0 2832 0 -1 770
box -8 -3 32 105
use NOR2X1  NOR2X1_148
timestamp 1711653199
transform 1 0 2672 0 -1 1170
box -8 -3 32 105
use NOR2X1  NOR2X1_149
timestamp 1711653199
transform 1 0 2440 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_150
timestamp 1711653199
transform 1 0 2936 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_151
timestamp 1711653199
transform 1 0 2304 0 -1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_152
timestamp 1711653199
transform 1 0 2856 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_153
timestamp 1711653199
transform 1 0 2368 0 1 1970
box -8 -3 32 105
use NOR2X1  NOR2X1_154
timestamp 1711653199
transform 1 0 2520 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_155
timestamp 1711653199
transform 1 0 3080 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_156
timestamp 1711653199
transform 1 0 3224 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_157
timestamp 1711653199
transform 1 0 3344 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_158
timestamp 1711653199
transform 1 0 3360 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_159
timestamp 1711653199
transform 1 0 3144 0 1 2170
box -8 -3 32 105
use NOR2X1  NOR2X1_160
timestamp 1711653199
transform 1 0 2368 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_161
timestamp 1711653199
transform 1 0 2320 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_162
timestamp 1711653199
transform 1 0 2248 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_163
timestamp 1711653199
transform 1 0 1368 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_164
timestamp 1711653199
transform 1 0 2064 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_165
timestamp 1711653199
transform 1 0 1736 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_166
timestamp 1711653199
transform 1 0 1600 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_167
timestamp 1711653199
transform 1 0 1672 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_168
timestamp 1711653199
transform 1 0 1480 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_169
timestamp 1711653199
transform 1 0 1416 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_170
timestamp 1711653199
transform 1 0 1248 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_171
timestamp 1711653199
transform 1 0 1240 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_172
timestamp 1711653199
transform 1 0 1392 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_173
timestamp 1711653199
transform 1 0 632 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_174
timestamp 1711653199
transform 1 0 560 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_175
timestamp 1711653199
transform 1 0 496 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_176
timestamp 1711653199
transform 1 0 512 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_177
timestamp 1711653199
transform 1 0 1464 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_178
timestamp 1711653199
transform 1 0 1632 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_179
timestamp 1711653199
transform 1 0 1688 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_180
timestamp 1711653199
transform 1 0 1624 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_181
timestamp 1711653199
transform 1 0 1216 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_182
timestamp 1711653199
transform 1 0 1192 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_183
timestamp 1711653199
transform 1 0 1160 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_184
timestamp 1711653199
transform 1 0 1288 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_185
timestamp 1711653199
transform 1 0 1152 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_186
timestamp 1711653199
transform 1 0 1200 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_187
timestamp 1711653199
transform 1 0 1720 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_188
timestamp 1711653199
transform 1 0 1056 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_189
timestamp 1711653199
transform 1 0 1120 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_190
timestamp 1711653199
transform 1 0 1144 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_191
timestamp 1711653199
transform 1 0 768 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_192
timestamp 1711653199
transform 1 0 704 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_193
timestamp 1711653199
transform 1 0 1920 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_194
timestamp 1711653199
transform 1 0 3144 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_195
timestamp 1711653199
transform 1 0 2008 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_196
timestamp 1711653199
transform 1 0 1800 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_197
timestamp 1711653199
transform 1 0 1776 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_198
timestamp 1711653199
transform 1 0 1488 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_199
timestamp 1711653199
transform 1 0 936 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_200
timestamp 1711653199
transform 1 0 688 0 1 2370
box -8 -3 32 105
use NOR2X1  NOR2X1_201
timestamp 1711653199
transform 1 0 344 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_202
timestamp 1711653199
transform 1 0 512 0 -1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_203
timestamp 1711653199
transform 1 0 192 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_204
timestamp 1711653199
transform 1 0 200 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_205
timestamp 1711653199
transform 1 0 224 0 1 2570
box -8 -3 32 105
use NOR2X1  NOR2X1_206
timestamp 1711653199
transform 1 0 208 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_207
timestamp 1711653199
transform 1 0 240 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_208
timestamp 1711653199
transform 1 0 288 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_209
timestamp 1711653199
transform 1 0 384 0 1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_210
timestamp 1711653199
transform 1 0 760 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_211
timestamp 1711653199
transform 1 0 1112 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_212
timestamp 1711653199
transform 1 0 776 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_213
timestamp 1711653199
transform 1 0 952 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_214
timestamp 1711653199
transform 1 0 1280 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_215
timestamp 1711653199
transform 1 0 1496 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_216
timestamp 1711653199
transform 1 0 1728 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_217
timestamp 1711653199
transform 1 0 1616 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_218
timestamp 1711653199
transform 1 0 1856 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_219
timestamp 1711653199
transform 1 0 1928 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_220
timestamp 1711653199
transform 1 0 2280 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_221
timestamp 1711653199
transform 1 0 2128 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_222
timestamp 1711653199
transform 1 0 2304 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_223
timestamp 1711653199
transform 1 0 2408 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_224
timestamp 1711653199
transform 1 0 2024 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_225
timestamp 1711653199
transform 1 0 2840 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_226
timestamp 1711653199
transform 1 0 3040 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_227
timestamp 1711653199
transform 1 0 3264 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_228
timestamp 1711653199
transform 1 0 3240 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_229
timestamp 1711653199
transform 1 0 3288 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_230
timestamp 1711653199
transform 1 0 3176 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_231
timestamp 1711653199
transform 1 0 3200 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_232
timestamp 1711653199
transform 1 0 3136 0 -1 2970
box -8 -3 32 105
use NOR2X1  NOR2X1_233
timestamp 1711653199
transform 1 0 3312 0 1 2770
box -8 -3 32 105
use OAI21X1  OAI21X1_0
timestamp 1711653199
transform 1 0 2936 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_1
timestamp 1711653199
transform 1 0 1608 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_2
timestamp 1711653199
transform 1 0 2456 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_3
timestamp 1711653199
transform 1 0 2272 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_4
timestamp 1711653199
transform 1 0 2136 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_5
timestamp 1711653199
transform 1 0 2760 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_6
timestamp 1711653199
transform 1 0 3072 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_7
timestamp 1711653199
transform 1 0 1160 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_8
timestamp 1711653199
transform 1 0 976 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_9
timestamp 1711653199
transform 1 0 560 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_10
timestamp 1711653199
transform 1 0 616 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_11
timestamp 1711653199
transform 1 0 2624 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_12
timestamp 1711653199
transform 1 0 544 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_13
timestamp 1711653199
transform 1 0 560 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_14
timestamp 1711653199
transform 1 0 1024 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_15
timestamp 1711653199
transform 1 0 1024 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_16
timestamp 1711653199
transform 1 0 2944 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_17
timestamp 1711653199
transform 1 0 1712 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_18
timestamp 1711653199
transform 1 0 2776 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_19
timestamp 1711653199
transform 1 0 736 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_20
timestamp 1711653199
transform 1 0 744 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_21
timestamp 1711653199
transform 1 0 2000 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_22
timestamp 1711653199
transform 1 0 1776 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_23
timestamp 1711653199
transform 1 0 1448 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_24
timestamp 1711653199
transform 1 0 1080 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_25
timestamp 1711653199
transform 1 0 1320 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_26
timestamp 1711653199
transform 1 0 2008 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_27
timestamp 1711653199
transform 1 0 1792 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_28
timestamp 1711653199
transform 1 0 232 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_29
timestamp 1711653199
transform 1 0 2200 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_30
timestamp 1711653199
transform 1 0 3032 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_31
timestamp 1711653199
transform 1 0 1432 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_32
timestamp 1711653199
transform 1 0 1472 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_33
timestamp 1711653199
transform 1 0 2632 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_34
timestamp 1711653199
transform 1 0 712 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_35
timestamp 1711653199
transform 1 0 672 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_36
timestamp 1711653199
transform 1 0 1072 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_37
timestamp 1711653199
transform 1 0 1080 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_38
timestamp 1711653199
transform 1 0 3072 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_39
timestamp 1711653199
transform 1 0 2464 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_40
timestamp 1711653199
transform 1 0 2488 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_41
timestamp 1711653199
transform 1 0 1376 0 -1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1711653199
transform 1 0 1480 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_43
timestamp 1711653199
transform 1 0 2336 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_44
timestamp 1711653199
transform 1 0 3056 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_45
timestamp 1711653199
transform 1 0 992 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_46
timestamp 1711653199
transform 1 0 1336 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_47
timestamp 1711653199
transform 1 0 2008 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_48
timestamp 1711653199
transform 1 0 1840 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_49
timestamp 1711653199
transform 1 0 1536 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_50
timestamp 1711653199
transform 1 0 1896 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_51
timestamp 1711653199
transform 1 0 1464 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_52
timestamp 1711653199
transform 1 0 2528 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_53
timestamp 1711653199
transform 1 0 1896 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_54
timestamp 1711653199
transform 1 0 496 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_55
timestamp 1711653199
transform 1 0 472 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_56
timestamp 1711653199
transform 1 0 2944 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_57
timestamp 1711653199
transform 1 0 792 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_58
timestamp 1711653199
transform 1 0 816 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_59
timestamp 1711653199
transform 1 0 1456 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_60
timestamp 1711653199
transform 1 0 824 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_61
timestamp 1711653199
transform 1 0 1536 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_62
timestamp 1711653199
transform 1 0 2072 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_63
timestamp 1711653199
transform 1 0 2568 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_64
timestamp 1711653199
transform 1 0 2008 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_65
timestamp 1711653199
transform 1 0 96 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_66
timestamp 1711653199
transform 1 0 1568 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_67
timestamp 1711653199
transform 1 0 3040 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_68
timestamp 1711653199
transform 1 0 1416 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_69
timestamp 1711653199
transform 1 0 1344 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_70
timestamp 1711653199
transform 1 0 2152 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_71
timestamp 1711653199
transform 1 0 2160 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_72
timestamp 1711653199
transform 1 0 2128 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_73
timestamp 1711653199
transform 1 0 2368 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_74
timestamp 1711653199
transform 1 0 2128 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_75
timestamp 1711653199
transform 1 0 1952 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_76
timestamp 1711653199
transform 1 0 2112 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_77
timestamp 1711653199
transform 1 0 2064 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_78
timestamp 1711653199
transform 1 0 2224 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_79
timestamp 1711653199
transform 1 0 2224 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_80
timestamp 1711653199
transform 1 0 2432 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_81
timestamp 1711653199
transform 1 0 2328 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_82
timestamp 1711653199
transform 1 0 2296 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_83
timestamp 1711653199
transform 1 0 2008 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_84
timestamp 1711653199
transform 1 0 2000 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_85
timestamp 1711653199
transform 1 0 2256 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_86
timestamp 1711653199
transform 1 0 2264 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_87
timestamp 1711653199
transform 1 0 2480 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_88
timestamp 1711653199
transform 1 0 2360 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_89
timestamp 1711653199
transform 1 0 2328 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_90
timestamp 1711653199
transform 1 0 2016 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_91
timestamp 1711653199
transform 1 0 1904 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_92
timestamp 1711653199
transform 1 0 2024 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_93
timestamp 1711653199
transform 1 0 1912 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_94
timestamp 1711653199
transform 1 0 2088 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_95
timestamp 1711653199
transform 1 0 2120 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_96
timestamp 1711653199
transform 1 0 1912 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_97
timestamp 1711653199
transform 1 0 1992 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_98
timestamp 1711653199
transform 1 0 2160 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_99
timestamp 1711653199
transform 1 0 1656 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_100
timestamp 1711653199
transform 1 0 1768 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_101
timestamp 1711653199
transform 1 0 1728 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_102
timestamp 1711653199
transform 1 0 2128 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_103
timestamp 1711653199
transform 1 0 2096 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_104
timestamp 1711653199
transform 1 0 1856 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_105
timestamp 1711653199
transform 1 0 1800 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_106
timestamp 1711653199
transform 1 0 1592 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_107
timestamp 1711653199
transform 1 0 1856 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_108
timestamp 1711653199
transform 1 0 1448 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_109
timestamp 1711653199
transform 1 0 1536 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_110
timestamp 1711653199
transform 1 0 1592 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_111
timestamp 1711653199
transform 1 0 1936 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_112
timestamp 1711653199
transform 1 0 2000 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_113
timestamp 1711653199
transform 1 0 1560 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_114
timestamp 1711653199
transform 1 0 1688 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_115
timestamp 1711653199
transform 1 0 1280 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_116
timestamp 1711653199
transform 1 0 1272 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_117
timestamp 1711653199
transform 1 0 1544 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_118
timestamp 1711653199
transform 1 0 1544 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_119
timestamp 1711653199
transform 1 0 1792 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_120
timestamp 1711653199
transform 1 0 1896 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_121
timestamp 1711653199
transform 1 0 1504 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_122
timestamp 1711653199
transform 1 0 1592 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_123
timestamp 1711653199
transform 1 0 1272 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_124
timestamp 1711653199
transform 1 0 1112 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_125
timestamp 1711653199
transform 1 0 2000 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_126
timestamp 1711653199
transform 1 0 2168 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_127
timestamp 1711653199
transform 1 0 2152 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_128
timestamp 1711653199
transform 1 0 1920 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_129
timestamp 1711653199
transform 1 0 1136 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_130
timestamp 1711653199
transform 1 0 1856 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_131
timestamp 1711653199
transform 1 0 336 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_132
timestamp 1711653199
transform 1 0 448 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_133
timestamp 1711653199
transform 1 0 640 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_134
timestamp 1711653199
transform 1 0 600 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_135
timestamp 1711653199
transform 1 0 672 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_136
timestamp 1711653199
transform 1 0 1008 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_137
timestamp 1711653199
transform 1 0 232 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_138
timestamp 1711653199
transform 1 0 96 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_139
timestamp 1711653199
transform 1 0 216 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_140
timestamp 1711653199
transform 1 0 168 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_141
timestamp 1711653199
transform 1 0 312 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_142
timestamp 1711653199
transform 1 0 528 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_143
timestamp 1711653199
transform 1 0 200 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_144
timestamp 1711653199
transform 1 0 80 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_145
timestamp 1711653199
transform 1 0 80 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_146
timestamp 1711653199
transform 1 0 104 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_147
timestamp 1711653199
transform 1 0 80 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_148
timestamp 1711653199
transform 1 0 96 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_149
timestamp 1711653199
transform 1 0 88 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_150
timestamp 1711653199
transform 1 0 448 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_151
timestamp 1711653199
transform 1 0 448 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_152
timestamp 1711653199
transform 1 0 392 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_153
timestamp 1711653199
transform 1 0 880 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_154
timestamp 1711653199
transform 1 0 480 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_155
timestamp 1711653199
transform 1 0 512 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_156
timestamp 1711653199
transform 1 0 680 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_157
timestamp 1711653199
transform 1 0 696 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_158
timestamp 1711653199
transform 1 0 816 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_159
timestamp 1711653199
transform 1 0 880 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_160
timestamp 1711653199
transform 1 0 1000 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_161
timestamp 1711653199
transform 1 0 616 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_162
timestamp 1711653199
transform 1 0 1072 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_163
timestamp 1711653199
transform 1 0 416 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_164
timestamp 1711653199
transform 1 0 408 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_165
timestamp 1711653199
transform 1 0 600 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_166
timestamp 1711653199
transform 1 0 488 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_167
timestamp 1711653199
transform 1 0 568 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_168
timestamp 1711653199
transform 1 0 808 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_169
timestamp 1711653199
transform 1 0 800 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_170
timestamp 1711653199
transform 1 0 608 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_171
timestamp 1711653199
transform 1 0 528 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_172
timestamp 1711653199
transform 1 0 488 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_173
timestamp 1711653199
transform 1 0 904 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_174
timestamp 1711653199
transform 1 0 568 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_175
timestamp 1711653199
transform 1 0 584 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_176
timestamp 1711653199
transform 1 0 864 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_177
timestamp 1711653199
transform 1 0 1000 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_178
timestamp 1711653199
transform 1 0 552 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_179
timestamp 1711653199
transform 1 0 952 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_180
timestamp 1711653199
transform 1 0 1736 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_181
timestamp 1711653199
transform 1 0 1728 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_182
timestamp 1711653199
transform 1 0 1000 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_183
timestamp 1711653199
transform 1 0 1656 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_184
timestamp 1711653199
transform 1 0 920 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_185
timestamp 1711653199
transform 1 0 888 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_186
timestamp 1711653199
transform 1 0 824 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_187
timestamp 1711653199
transform 1 0 752 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_188
timestamp 1711653199
transform 1 0 792 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_189
timestamp 1711653199
transform 1 0 928 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_190
timestamp 1711653199
transform 1 0 624 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_191
timestamp 1711653199
transform 1 0 456 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_192
timestamp 1711653199
transform 1 0 416 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_193
timestamp 1711653199
transform 1 0 400 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_194
timestamp 1711653199
transform 1 0 480 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_195
timestamp 1711653199
transform 1 0 712 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_196
timestamp 1711653199
transform 1 0 560 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_197
timestamp 1711653199
transform 1 0 136 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_198
timestamp 1711653199
transform 1 0 328 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_199
timestamp 1711653199
transform 1 0 296 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_200
timestamp 1711653199
transform 1 0 256 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_201
timestamp 1711653199
transform 1 0 592 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_202
timestamp 1711653199
transform 1 0 1416 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_203
timestamp 1711653199
transform 1 0 1392 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_204
timestamp 1711653199
transform 1 0 1368 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_205
timestamp 1711653199
transform 1 0 1448 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_206
timestamp 1711653199
transform 1 0 1456 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_207
timestamp 1711653199
transform 1 0 1424 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_208
timestamp 1711653199
transform 1 0 1312 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_209
timestamp 1711653199
transform 1 0 1144 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_210
timestamp 1711653199
transform 1 0 928 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_211
timestamp 1711653199
transform 1 0 1056 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_212
timestamp 1711653199
transform 1 0 952 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_213
timestamp 1711653199
transform 1 0 928 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_214
timestamp 1711653199
transform 1 0 1280 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_215
timestamp 1711653199
transform 1 0 1336 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_216
timestamp 1711653199
transform 1 0 1280 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_217
timestamp 1711653199
transform 1 0 1808 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_218
timestamp 1711653199
transform 1 0 1624 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_219
timestamp 1711653199
transform 1 0 1320 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_220
timestamp 1711653199
transform 1 0 1192 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_221
timestamp 1711653199
transform 1 0 1192 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_222
timestamp 1711653199
transform 1 0 1176 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_223
timestamp 1711653199
transform 1 0 1296 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_224
timestamp 1711653199
transform 1 0 1216 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_225
timestamp 1711653199
transform 1 0 1416 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_226
timestamp 1711653199
transform 1 0 1688 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_227
timestamp 1711653199
transform 1 0 1384 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_228
timestamp 1711653199
transform 1 0 1072 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_229
timestamp 1711653199
transform 1 0 1080 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_230
timestamp 1711653199
transform 1 0 1024 0 1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_231
timestamp 1711653199
transform 1 0 1064 0 1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_232
timestamp 1711653199
transform 1 0 1136 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_233
timestamp 1711653199
transform 1 0 1064 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_234
timestamp 1711653199
transform 1 0 1344 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_235
timestamp 1711653199
transform 1 0 1776 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_236
timestamp 1711653199
transform 1 0 2240 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_237
timestamp 1711653199
transform 1 0 2400 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_238
timestamp 1711653199
transform 1 0 2320 0 -1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_239
timestamp 1711653199
transform 1 0 2232 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_240
timestamp 1711653199
transform 1 0 2024 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_241
timestamp 1711653199
transform 1 0 2272 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_242
timestamp 1711653199
transform 1 0 2008 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_243
timestamp 1711653199
transform 1 0 2272 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_244
timestamp 1711653199
transform 1 0 3040 0 -1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_245
timestamp 1711653199
transform 1 0 3136 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_246
timestamp 1711653199
transform 1 0 3184 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_247
timestamp 1711653199
transform 1 0 3096 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_248
timestamp 1711653199
transform 1 0 2512 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_249
timestamp 1711653199
transform 1 0 2584 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_250
timestamp 1711653199
transform 1 0 3272 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_251
timestamp 1711653199
transform 1 0 3288 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_252
timestamp 1711653199
transform 1 0 3296 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_253
timestamp 1711653199
transform 1 0 3216 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_254
timestamp 1711653199
transform 1 0 2928 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_255
timestamp 1711653199
transform 1 0 2648 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_256
timestamp 1711653199
transform 1 0 3144 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_257
timestamp 1711653199
transform 1 0 3352 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_258
timestamp 1711653199
transform 1 0 3352 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_259
timestamp 1711653199
transform 1 0 3352 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_260
timestamp 1711653199
transform 1 0 2832 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_261
timestamp 1711653199
transform 1 0 2400 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_262
timestamp 1711653199
transform 1 0 2704 0 1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_263
timestamp 1711653199
transform 1 0 2656 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_264
timestamp 1711653199
transform 1 0 2824 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_265
timestamp 1711653199
transform 1 0 2704 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_266
timestamp 1711653199
transform 1 0 2720 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_267
timestamp 1711653199
transform 1 0 2736 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_268
timestamp 1711653199
transform 1 0 2560 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_269
timestamp 1711653199
transform 1 0 2784 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_270
timestamp 1711653199
transform 1 0 2320 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_271
timestamp 1711653199
transform 1 0 2704 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_272
timestamp 1711653199
transform 1 0 2688 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_273
timestamp 1711653199
transform 1 0 2736 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_274
timestamp 1711653199
transform 1 0 2744 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_275
timestamp 1711653199
transform 1 0 2712 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_276
timestamp 1711653199
transform 1 0 2672 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_277
timestamp 1711653199
transform 1 0 2672 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_278
timestamp 1711653199
transform 1 0 2640 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_279
timestamp 1711653199
transform 1 0 2328 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_280
timestamp 1711653199
transform 1 0 2360 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_281
timestamp 1711653199
transform 1 0 2448 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_282
timestamp 1711653199
transform 1 0 2912 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_283
timestamp 1711653199
transform 1 0 2832 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_284
timestamp 1711653199
transform 1 0 2904 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_285
timestamp 1711653199
transform 1 0 2664 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_286
timestamp 1711653199
transform 1 0 2568 0 -1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_287
timestamp 1711653199
transform 1 0 2632 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_288
timestamp 1711653199
transform 1 0 2456 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_289
timestamp 1711653199
transform 1 0 2424 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_290
timestamp 1711653199
transform 1 0 2440 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_291
timestamp 1711653199
transform 1 0 2888 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_292
timestamp 1711653199
transform 1 0 2856 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_293
timestamp 1711653199
transform 1 0 2912 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_294
timestamp 1711653199
transform 1 0 2864 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_295
timestamp 1711653199
transform 1 0 2800 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_296
timestamp 1711653199
transform 1 0 2728 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_297
timestamp 1711653199
transform 1 0 2824 0 1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_298
timestamp 1711653199
transform 1 0 2664 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_299
timestamp 1711653199
transform 1 0 2360 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_300
timestamp 1711653199
transform 1 0 2408 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_301
timestamp 1711653199
transform 1 0 3072 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_302
timestamp 1711653199
transform 1 0 3000 0 -1 1570
box -8 -3 34 105
use OAI21X1  OAI21X1_303
timestamp 1711653199
transform 1 0 3000 0 -1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_304
timestamp 1711653199
transform 1 0 3016 0 1 970
box -8 -3 34 105
use OAI21X1  OAI21X1_305
timestamp 1711653199
transform 1 0 2984 0 1 1170
box -8 -3 34 105
use OAI21X1  OAI21X1_306
timestamp 1711653199
transform 1 0 3056 0 1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_307
timestamp 1711653199
transform 1 0 3080 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_308
timestamp 1711653199
transform 1 0 2992 0 1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_309
timestamp 1711653199
transform 1 0 3024 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_310
timestamp 1711653199
transform 1 0 2760 0 -1 1970
box -8 -3 34 105
use OAI21X1  OAI21X1_311
timestamp 1711653199
transform 1 0 2936 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_312
timestamp 1711653199
transform 1 0 2928 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_313
timestamp 1711653199
transform 1 0 3144 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_314
timestamp 1711653199
transform 1 0 3104 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_315
timestamp 1711653199
transform 1 0 3064 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_316
timestamp 1711653199
transform 1 0 3296 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_317
timestamp 1711653199
transform 1 0 3328 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_318
timestamp 1711653199
transform 1 0 2704 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_319
timestamp 1711653199
transform 1 0 2736 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_320
timestamp 1711653199
transform 1 0 2904 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_321
timestamp 1711653199
transform 1 0 3104 0 1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_322
timestamp 1711653199
transform 1 0 3136 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_323
timestamp 1711653199
transform 1 0 3208 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_324
timestamp 1711653199
transform 1 0 3136 0 -1 2370
box -8 -3 34 105
use OAI21X1  OAI21X1_325
timestamp 1711653199
transform 1 0 3192 0 1 2170
box -8 -3 34 105
use OAI21X1  OAI21X1_326
timestamp 1711653199
transform 1 0 2624 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_327
timestamp 1711653199
transform 1 0 2640 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_328
timestamp 1711653199
transform 1 0 2032 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_329
timestamp 1711653199
transform 1 0 2376 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_330
timestamp 1711653199
transform 1 0 2480 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_331
timestamp 1711653199
transform 1 0 2160 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_332
timestamp 1711653199
transform 1 0 1392 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_333
timestamp 1711653199
transform 1 0 1432 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_334
timestamp 1711653199
transform 1 0 1656 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_335
timestamp 1711653199
transform 1 0 1816 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_336
timestamp 1711653199
transform 1 0 1784 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_337
timestamp 1711653199
transform 1 0 1584 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_338
timestamp 1711653199
transform 1 0 1624 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_339
timestamp 1711653199
transform 1 0 1696 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_340
timestamp 1711653199
transform 1 0 1696 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_341
timestamp 1711653199
transform 1 0 1464 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_342
timestamp 1711653199
transform 1 0 1536 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_343
timestamp 1711653199
transform 1 0 1400 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_344
timestamp 1711653199
transform 1 0 1368 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_345
timestamp 1711653199
transform 1 0 1304 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_346
timestamp 1711653199
transform 1 0 1344 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_347
timestamp 1711653199
transform 1 0 1040 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_348
timestamp 1711653199
transform 1 0 1072 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_349
timestamp 1711653199
transform 1 0 920 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_350
timestamp 1711653199
transform 1 0 976 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_351
timestamp 1711653199
transform 1 0 1160 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_352
timestamp 1711653199
transform 1 0 1192 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_353
timestamp 1711653199
transform 1 0 696 0 1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_354
timestamp 1711653199
transform 1 0 632 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_355
timestamp 1711653199
transform 1 0 488 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_356
timestamp 1711653199
transform 1 0 552 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_357
timestamp 1711653199
transform 1 0 328 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_358
timestamp 1711653199
transform 1 0 528 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_359
timestamp 1711653199
transform 1 0 248 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_360
timestamp 1711653199
transform 1 0 560 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_361
timestamp 1711653199
transform 1 0 864 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_362
timestamp 1711653199
transform 1 0 800 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_363
timestamp 1711653199
transform 1 0 200 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_364
timestamp 1711653199
transform 1 0 600 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_365
timestamp 1711653199
transform 1 0 408 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_366
timestamp 1711653199
transform 1 0 528 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_367
timestamp 1711653199
transform 1 0 216 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_368
timestamp 1711653199
transform 1 0 440 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_369
timestamp 1711653199
transform 1 0 216 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_370
timestamp 1711653199
transform 1 0 480 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_371
timestamp 1711653199
transform 1 0 528 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_372
timestamp 1711653199
transform 1 0 672 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_373
timestamp 1711653199
transform 1 0 360 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_374
timestamp 1711653199
transform 1 0 640 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_375
timestamp 1711653199
transform 1 0 688 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_376
timestamp 1711653199
transform 1 0 720 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_377
timestamp 1711653199
transform 1 0 904 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_378
timestamp 1711653199
transform 1 0 888 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_379
timestamp 1711653199
transform 1 0 1032 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_380
timestamp 1711653199
transform 1 0 1064 0 -1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_381
timestamp 1711653199
transform 1 0 1384 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_382
timestamp 1711653199
transform 1 0 1424 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_383
timestamp 1711653199
transform 1 0 1560 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_384
timestamp 1711653199
transform 1 0 1528 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_385
timestamp 1711653199
transform 1 0 1744 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_386
timestamp 1711653199
transform 1 0 1656 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_387
timestamp 1711653199
transform 1 0 1832 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_388
timestamp 1711653199
transform 1 0 1648 0 1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_389
timestamp 1711653199
transform 1 0 2976 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_390
timestamp 1711653199
transform 1 0 3008 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_391
timestamp 1711653199
transform 1 0 3184 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_392
timestamp 1711653199
transform 1 0 3216 0 1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_393
timestamp 1711653199
transform 1 0 3264 0 -1 3170
box -8 -3 34 105
use OAI21X1  OAI21X1_394
timestamp 1711653199
transform 1 0 3088 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_395
timestamp 1711653199
transform 1 0 2976 0 1 2770
box -8 -3 34 105
use OAI22X1  OAI22X1_0
timestamp 1711653199
transform 1 0 2416 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_1
timestamp 1711653199
transform 1 0 2200 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_2
timestamp 1711653199
transform 1 0 2520 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_3
timestamp 1711653199
transform 1 0 2496 0 -1 1370
box -8 -3 46 105
use OAI22X1  OAI22X1_4
timestamp 1711653199
transform 1 0 2048 0 -1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_5
timestamp 1711653199
transform 1 0 2000 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_6
timestamp 1711653199
transform 1 0 1824 0 1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_7
timestamp 1711653199
transform 1 0 968 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_8
timestamp 1711653199
transform 1 0 672 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_9
timestamp 1711653199
transform 1 0 736 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_10
timestamp 1711653199
transform 1 0 800 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_11
timestamp 1711653199
transform 1 0 936 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_12
timestamp 1711653199
transform 1 0 816 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_13
timestamp 1711653199
transform 1 0 704 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_14
timestamp 1711653199
transform 1 0 752 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_15
timestamp 1711653199
transform 1 0 1528 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_16
timestamp 1711653199
transform 1 0 752 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_17
timestamp 1711653199
transform 1 0 648 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_18
timestamp 1711653199
transform 1 0 648 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_19
timestamp 1711653199
transform 1 0 1368 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_20
timestamp 1711653199
transform 1 0 1168 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_21
timestamp 1711653199
transform 1 0 1232 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_22
timestamp 1711653199
transform 1 0 1272 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_23
timestamp 1711653199
transform 1 0 1768 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_24
timestamp 1711653199
transform 1 0 936 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_25
timestamp 1711653199
transform 1 0 1856 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_26
timestamp 1711653199
transform 1 0 2112 0 -1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_27
timestamp 1711653199
transform 1 0 2216 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_28
timestamp 1711653199
transform 1 0 3120 0 1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_29
timestamp 1711653199
transform 1 0 2440 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_30
timestamp 1711653199
transform 1 0 2352 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_31
timestamp 1711653199
transform 1 0 2824 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_32
timestamp 1711653199
transform 1 0 2800 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_33
timestamp 1711653199
transform 1 0 2856 0 -1 1770
box -8 -3 46 105
use OAI22X1  OAI22X1_34
timestamp 1711653199
transform 1 0 2616 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_35
timestamp 1711653199
transform 1 0 1744 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_36
timestamp 1711653199
transform 1 0 2536 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_37
timestamp 1711653199
transform 1 0 1696 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_38
timestamp 1711653199
transform 1 0 2840 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_39
timestamp 1711653199
transform 1 0 1192 0 -1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_40
timestamp 1711653199
transform 1 0 3088 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_41
timestamp 1711653199
transform 1 0 3128 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_42
timestamp 1711653199
transform 1 0 2808 0 1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_43
timestamp 1711653199
transform 1 0 2792 0 -1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_44
timestamp 1711653199
transform 1 0 3320 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_45
timestamp 1711653199
transform 1 0 3264 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_46
timestamp 1711653199
transform 1 0 3240 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_47
timestamp 1711653199
transform 1 0 3192 0 1 2370
box -8 -3 46 105
use OAI22X1  OAI22X1_48
timestamp 1711653199
transform 1 0 2208 0 -1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_49
timestamp 1711653199
transform 1 0 1160 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_50
timestamp 1711653199
transform 1 0 1952 0 -1 3170
box -8 -3 46 105
use OAI22X1  OAI22X1_51
timestamp 1711653199
transform 1 0 1864 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_52
timestamp 1711653199
transform 1 0 1760 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_53
timestamp 1711653199
transform 1 0 1824 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_54
timestamp 1711653199
transform 1 0 1544 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_55
timestamp 1711653199
transform 1 0 1288 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_56
timestamp 1711653199
transform 1 0 1048 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_57
timestamp 1711653199
transform 1 0 960 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_58
timestamp 1711653199
transform 1 0 1192 0 1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_59
timestamp 1711653199
transform 1 0 656 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_60
timestamp 1711653199
transform 1 0 616 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_61
timestamp 1711653199
transform 1 0 656 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_62
timestamp 1711653199
transform 1 0 720 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_63
timestamp 1711653199
transform 1 0 1040 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_64
timestamp 1711653199
transform 1 0 1088 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_65
timestamp 1711653199
transform 1 0 1192 0 -1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_66
timestamp 1711653199
transform 1 0 1264 0 1 2570
box -8 -3 46 105
use OAI22X1  OAI22X1_67
timestamp 1711653199
transform 1 0 3248 0 1 2970
box -8 -3 46 105
use OR2X1  OR2X1_0
timestamp 1711653199
transform 1 0 3056 0 -1 1570
box -8 -3 40 105
use OR2X1  OR2X1_1
timestamp 1711653199
transform 1 0 3280 0 1 1770
box -8 -3 40 105
use OR2X1  OR2X1_2
timestamp 1711653199
transform 1 0 3208 0 1 1770
box -8 -3 40 105
use OR2X1  OR2X1_3
timestamp 1711653199
transform 1 0 2816 0 -1 2170
box -8 -3 40 105
use OR2X1  OR2X1_4
timestamp 1711653199
transform 1 0 2728 0 -1 3170
box -8 -3 40 105
use OR2X1  OR2X1_5
timestamp 1711653199
transform 1 0 3128 0 1 1570
box -8 -3 40 105
use OR2X1  OR2X1_6
timestamp 1711653199
transform 1 0 2984 0 1 2370
box -8 -3 40 105
use OR2X1  OR2X1_7
timestamp 1711653199
transform 1 0 2848 0 1 970
box -8 -3 40 105
use OR2X1  OR2X1_8
timestamp 1711653199
transform 1 0 1464 0 1 1170
box -8 -3 40 105
use OR2X1  OR2X1_9
timestamp 1711653199
transform 1 0 2376 0 1 1170
box -8 -3 40 105
use OR2X1  OR2X1_10
timestamp 1711653199
transform 1 0 1960 0 -1 1770
box -8 -3 40 105
use OR2X1  OR2X1_11
timestamp 1711653199
transform 1 0 2048 0 -1 1770
box -8 -3 40 105
use OR2X1  OR2X1_12
timestamp 1711653199
transform 1 0 1992 0 -1 970
box -8 -3 40 105
use OR2X1  OR2X1_13
timestamp 1711653199
transform 1 0 2136 0 1 570
box -8 -3 40 105
use OR2X1  OR2X1_14
timestamp 1711653199
transform 1 0 2000 0 1 370
box -8 -3 40 105
use OR2X1  OR2X1_15
timestamp 1711653199
transform 1 0 352 0 1 770
box -8 -3 40 105
use OR2X1  OR2X1_16
timestamp 1711653199
transform 1 0 728 0 -1 570
box -8 -3 40 105
use OR2X1  OR2X1_17
timestamp 1711653199
transform 1 0 440 0 1 770
box -8 -3 40 105
use OR2X1  OR2X1_18
timestamp 1711653199
transform 1 0 600 0 -1 770
box -8 -3 40 105
use OR2X1  OR2X1_19
timestamp 1711653199
transform 1 0 848 0 1 970
box -8 -3 40 105
use OR2X1  OR2X1_20
timestamp 1711653199
transform 1 0 808 0 1 370
box -8 -3 40 105
use OR2X1  OR2X1_21
timestamp 1711653199
transform 1 0 144 0 -1 1170
box -8 -3 40 105
use OR2X1  OR2X1_22
timestamp 1711653199
transform 1 0 200 0 -1 1170
box -8 -3 40 105
use OR2X1  OR2X1_23
timestamp 1711653199
transform 1 0 1112 0 1 370
box -8 -3 40 105
use OR2X1  OR2X1_24
timestamp 1711653199
transform 1 0 1320 0 -1 570
box -8 -3 40 105
use OR2X1  OR2X1_25
timestamp 1711653199
transform 1 0 1056 0 -1 770
box -8 -3 40 105
use OR2X1  OR2X1_26
timestamp 1711653199
transform 1 0 2368 0 -1 170
box -8 -3 40 105
use OR2X1  OR2X1_27
timestamp 1711653199
transform 1 0 1928 0 1 2170
box -8 -3 40 105
use OR2X1  OR2X1_28
timestamp 1711653199
transform 1 0 3128 0 -1 570
box -8 -3 40 105
use OR2X1  OR2X1_29
timestamp 1711653199
transform 1 0 2736 0 1 170
box -8 -3 40 105
use OR2X1  OR2X1_30
timestamp 1711653199
transform 1 0 2408 0 -1 2170
box -8 -3 40 105
use OR2X1  OR2X1_31
timestamp 1711653199
transform 1 0 3264 0 1 2370
box -8 -3 40 105
use OR2X1  OR2X1_32
timestamp 1711653199
transform 1 0 1288 0 -1 2770
box -8 -3 40 105
use OR2X1  OR2X1_33
timestamp 1711653199
transform 1 0 3184 0 -1 3170
box -8 -3 40 105
use OR2X1  OR2X1_34
timestamp 1711653199
transform 1 0 3328 0 -1 3170
box -8 -3 40 105
use OR2X1  OR2X1_35
timestamp 1711653199
transform 1 0 3248 0 -1 2770
box -8 -3 40 105
use OR2X2  OR2X2_0
timestamp 1711653199
transform 1 0 3360 0 1 2770
box -7 -3 35 105
use OR2X2  OR2X2_1
timestamp 1711653199
transform 1 0 2608 0 -1 970
box -7 -3 35 105
use top_module_VIA0  top_module_VIA0_0
timestamp 1711653199
transform 1 0 3448 0 1 3317
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_1
timestamp 1711653199
transform 1 0 3448 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_2
timestamp 1711653199
transform 1 0 24 0 1 3317
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_3
timestamp 1711653199
transform 1 0 24 0 1 23
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_4
timestamp 1711653199
transform 1 0 3424 0 1 3293
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_5
timestamp 1711653199
transform 1 0 3424 0 1 47
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_6
timestamp 1711653199
transform 1 0 48 0 1 3293
box -10 -10 10 10
use top_module_VIA0  top_module_VIA0_7
timestamp 1711653199
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_module_VIA1  top_module_VIA1_0
timestamp 1711653199
transform 1 0 3448 0 1 3270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_1
timestamp 1711653199
transform 1 0 3448 0 1 3070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_2
timestamp 1711653199
transform 1 0 3448 0 1 2870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_3
timestamp 1711653199
transform 1 0 3448 0 1 2670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_4
timestamp 1711653199
transform 1 0 3448 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_5
timestamp 1711653199
transform 1 0 3448 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_6
timestamp 1711653199
transform 1 0 3448 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_7
timestamp 1711653199
transform 1 0 3448 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_8
timestamp 1711653199
transform 1 0 3448 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_9
timestamp 1711653199
transform 1 0 3448 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_10
timestamp 1711653199
transform 1 0 3448 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_11
timestamp 1711653199
transform 1 0 3448 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_12
timestamp 1711653199
transform 1 0 3448 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_13
timestamp 1711653199
transform 1 0 3448 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_14
timestamp 1711653199
transform 1 0 3448 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_15
timestamp 1711653199
transform 1 0 3448 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_16
timestamp 1711653199
transform 1 0 3448 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_17
timestamp 1711653199
transform 1 0 24 0 1 3270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_18
timestamp 1711653199
transform 1 0 24 0 1 3070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_19
timestamp 1711653199
transform 1 0 24 0 1 2870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_20
timestamp 1711653199
transform 1 0 24 0 1 2670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_21
timestamp 1711653199
transform 1 0 24 0 1 2470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_22
timestamp 1711653199
transform 1 0 24 0 1 2270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_23
timestamp 1711653199
transform 1 0 24 0 1 2070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_24
timestamp 1711653199
transform 1 0 24 0 1 1870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_25
timestamp 1711653199
transform 1 0 24 0 1 1670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_26
timestamp 1711653199
transform 1 0 24 0 1 1470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_27
timestamp 1711653199
transform 1 0 24 0 1 1270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_28
timestamp 1711653199
transform 1 0 24 0 1 1070
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_29
timestamp 1711653199
transform 1 0 24 0 1 870
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_30
timestamp 1711653199
transform 1 0 24 0 1 670
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_31
timestamp 1711653199
transform 1 0 24 0 1 470
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_32
timestamp 1711653199
transform 1 0 24 0 1 270
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_33
timestamp 1711653199
transform 1 0 24 0 1 70
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_34
timestamp 1711653199
transform 1 0 48 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_35
timestamp 1711653199
transform 1 0 48 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_36
timestamp 1711653199
transform 1 0 48 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_37
timestamp 1711653199
transform 1 0 48 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_38
timestamp 1711653199
transform 1 0 48 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_39
timestamp 1711653199
transform 1 0 48 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_40
timestamp 1711653199
transform 1 0 48 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_41
timestamp 1711653199
transform 1 0 48 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_42
timestamp 1711653199
transform 1 0 48 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_43
timestamp 1711653199
transform 1 0 48 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_44
timestamp 1711653199
transform 1 0 48 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_45
timestamp 1711653199
transform 1 0 48 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_46
timestamp 1711653199
transform 1 0 48 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_47
timestamp 1711653199
transform 1 0 48 0 1 2770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_48
timestamp 1711653199
transform 1 0 48 0 1 2970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_49
timestamp 1711653199
transform 1 0 48 0 1 3170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_50
timestamp 1711653199
transform 1 0 3424 0 1 170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_51
timestamp 1711653199
transform 1 0 3424 0 1 370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_52
timestamp 1711653199
transform 1 0 3424 0 1 570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_53
timestamp 1711653199
transform 1 0 3424 0 1 770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_54
timestamp 1711653199
transform 1 0 3424 0 1 970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_55
timestamp 1711653199
transform 1 0 3424 0 1 1170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_56
timestamp 1711653199
transform 1 0 3424 0 1 1370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_57
timestamp 1711653199
transform 1 0 3424 0 1 1570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_58
timestamp 1711653199
transform 1 0 3424 0 1 1770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_59
timestamp 1711653199
transform 1 0 3424 0 1 1970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_60
timestamp 1711653199
transform 1 0 3424 0 1 2170
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_61
timestamp 1711653199
transform 1 0 3424 0 1 2370
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_62
timestamp 1711653199
transform 1 0 3424 0 1 2570
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_63
timestamp 1711653199
transform 1 0 3424 0 1 2770
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_64
timestamp 1711653199
transform 1 0 3424 0 1 2970
box -10 -3 10 3
use top_module_VIA1  top_module_VIA1_65
timestamp 1711653199
transform 1 0 3424 0 1 3170
box -10 -3 10 3
use XNOR2X1  XNOR2X1_0
timestamp 1711653199
transform 1 0 2784 0 1 2570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_1
timestamp 1711653199
transform 1 0 2648 0 1 2170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_2
timestamp 1711653199
transform 1 0 2752 0 1 2170
box -8 -3 64 105
use XOR2X1  XOR2X1_0
timestamp 1711653199
transform 1 0 2680 0 -1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_1
timestamp 1711653199
transform 1 0 2648 0 1 2570
box -8 -3 64 105
use XOR2X1  XOR2X1_2
timestamp 1711653199
transform 1 0 2720 0 1 2970
box -8 -3 64 105
<< labels >>
rlabel metal1 2708 2935 2708 2935 4 in_clka
rlabel electrodecontact s 1788 2725 1788 2725 4 in_clkb
rlabel electrodecontact s 2468 3135 2468 3135 4 in_restart
rlabel electrodecontact s 3276 2805 3276 2805 4 in_move[1]
rlabel electrodecontact s 3348 2805 3348 2805 4 in_move[0]
rlabel metal1 1660 2415 1660 2415 4 board_out[31]
rlabel metal1 1716 2415 1716 2415 4 board_out[30]
rlabel electrodecontact s 1980 2325 1980 2325 4 board_out[29]
rlabel electrodecontact s 1740 2325 1740 2325 4 board_out[28]
rlabel metal1 1316 2615 1316 2615 4 board_out[27]
rlabel electrodecontact s 1188 2525 1188 2525 4 board_out[26]
rlabel metal1 1004 2525 1004 2525 4 board_out[25]
rlabel electrodecontact s 1020 2525 1020 2525 4 board_out[24]
rlabel metal1 1140 2615 1140 2615 4 board_out[23]
rlabel metal1 1156 2615 1156 2615 4 board_out[22]
rlabel electrodecontact s 276 2215 276 2215 4 board_out[21]
rlabel electrodecontact s 92 2125 92 2125 4 board_out[20]
rlabel electrodecontact s 764 2725 764 2725 4 board_out[19]
rlabel metal1 748 2725 748 2725 4 board_out[18]
rlabel metal1 764 2615 764 2615 4 board_out[17]
rlabel electrodecontact s 996 2615 996 2615 4 board_out[16]
rlabel metal1 772 2925 772 2925 4 board_out[15]
rlabel metal1 692 2925 692 2925 4 board_out[14]
rlabel metal1 828 3015 828 3015 4 board_out[13]
rlabel metal1 892 3015 892 3015 4 board_out[12]
rlabel electrodecontact s 948 3015 948 3015 4 board_out[11]
rlabel metal1 932 3015 932 3015 4 board_out[10]
rlabel metal1 1108 3015 1108 3015 4 board_out[9]
rlabel metal1 1244 3015 1244 3015 4 board_out[8]
rlabel metal1 1908 2925 1908 2925 4 board_out[7]
rlabel electrodecontact s 2164 2925 2164 2925 4 board_out[6]
rlabel electrodecontact s 2684 2925 2684 2925 4 board_out[5]
rlabel metal1 2140 3015 2140 3015 4 board_out[4]
rlabel electrodecontact s 2060 2925 2060 2925 4 board_out[3]
rlabel metal1 2572 3015 2572 3015 4 board_out[2]
rlabel metal1 2148 2925 2148 2925 4 board_out[1]
rlabel metal1 2076 3015 2076 3015 4 board_out[0]
rlabel metal2 38 37 38 37 4 gnd
rlabel metal2 14 13 14 13 4 vdd
<< properties >>
string path 26604.002 24435.000 26676.002 24435.000 
<< end >>
