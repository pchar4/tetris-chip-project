magic
tech scmos
timestamp 1710841341
<< nwell >>
rect -8 48 40 105
<< ntransistor >>
rect 7 6 9 26
rect 12 6 14 26
rect 20 6 22 26
<< ptransistor >>
rect 7 74 9 94
rect 15 74 17 94
rect 23 54 25 94
<< ndiffusion >>
rect 2 25 7 26
rect 6 6 7 25
rect 9 6 12 26
rect 14 25 20 26
rect 14 6 15 25
rect 19 6 20 25
rect 22 25 27 26
rect 22 6 23 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 74 7 93
rect 9 93 15 94
rect 9 74 10 93
rect 14 74 15 93
rect 17 92 23 94
rect 17 74 18 92
rect 22 58 23 92
rect 18 56 23 58
rect 20 54 23 56
rect 25 93 30 94
rect 25 54 26 93
<< ndcontact >>
rect 2 6 6 25
rect 15 6 19 25
rect 23 6 27 25
<< pdcontact >>
rect 2 74 6 93
rect 10 74 14 93
rect 18 58 22 92
rect 26 54 30 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 7 73 9 74
rect 5 71 9 73
rect 5 41 7 71
rect 6 37 7 41
rect 15 39 17 74
rect 5 30 7 37
rect 16 37 17 39
rect 5 28 9 30
rect 7 26 9 28
rect 12 26 14 35
rect 23 33 25 54
rect 24 31 25 33
rect 20 26 22 29
rect 7 4 9 6
rect 12 4 14 6
rect 20 4 22 6
<< polycontact >>
rect 2 37 6 41
rect 12 35 16 39
rect 20 29 24 33
<< metal1 >>
rect -2 102 34 103
rect 2 98 14 102
rect 18 98 34 102
rect -2 97 34 98
rect 2 93 6 97
rect 10 93 14 94
rect 11 53 14 74
rect 18 92 22 97
rect 18 56 22 58
rect 26 93 30 94
rect 11 50 23 53
rect 10 43 14 47
rect 2 33 6 37
rect 11 39 14 43
rect 11 36 12 39
rect 20 33 23 50
rect 27 47 30 54
rect 26 43 30 47
rect 9 30 20 32
rect 3 29 20 30
rect 3 27 12 29
rect 3 26 6 27
rect 27 26 30 43
rect 2 25 6 26
rect 23 25 30 26
rect 27 21 30 25
rect 15 3 19 6
rect -2 2 34 3
rect 2 -2 14 2
rect 18 -2 34 2
rect -2 -3 34 -2
<< m1p >>
rect 10 43 14 47
rect 26 43 30 47
rect 2 33 6 37
<< labels >>
rlabel metal1 4 100 4 100 4 vdd
rlabel metal1 4 0 4 0 4 gnd
rlabel metal1 4 35 4 35 4 A
rlabel metal1 12 45 12 45 4 B
rlabel metal1 28 45 28 45 4 Y
<< end >>
