magic
tech scmos
timestamp 1710841341
<< nwell >>
rect -7 48 39 105
<< ntransistor >>
rect 10 6 12 26
rect 15 6 17 26
rect 23 6 25 16
<< ptransistor >>
rect 7 54 9 94
rect 15 54 17 94
rect 23 54 25 94
<< ndiffusion >>
rect 5 25 10 26
rect 9 6 10 25
rect 12 6 15 26
rect 17 25 22 26
rect 17 6 18 25
rect 22 6 23 16
rect 25 15 30 16
rect 25 6 26 15
<< pdiffusion >>
rect 2 92 7 94
rect 6 58 7 92
rect 2 54 7 58
rect 9 60 10 94
rect 14 60 15 94
rect 9 54 15 60
rect 17 93 23 94
rect 17 54 18 93
rect 22 54 23 93
rect 25 93 30 94
rect 25 54 26 93
<< ndcontact >>
rect 5 6 9 25
rect 18 6 22 25
rect 26 6 30 15
<< pdcontact >>
rect 2 58 6 92
rect 10 60 14 94
rect 18 54 22 93
rect 26 54 30 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 7 49 9 54
rect 4 29 6 47
rect 15 41 17 54
rect 14 37 17 41
rect 4 27 12 29
rect 10 26 12 27
rect 15 26 17 37
rect 23 16 25 54
rect 10 4 12 6
rect 15 4 17 6
rect 23 4 25 6
<< polycontact >>
rect 6 45 10 49
rect 10 37 14 41
rect 25 19 29 23
<< metal1 >>
rect -2 102 34 103
rect 2 98 14 102
rect 18 98 34 102
rect -2 97 34 98
rect 10 94 14 97
rect 2 92 6 94
rect 18 93 22 94
rect 2 57 6 58
rect 2 54 18 57
rect 26 93 30 94
rect 2 45 6 47
rect 26 47 29 54
rect 2 44 10 45
rect 18 44 30 47
rect 2 43 6 44
rect 10 33 14 37
rect 18 26 21 44
rect 26 43 30 44
rect 5 25 9 26
rect 18 25 22 26
rect 26 23 30 27
rect 26 15 30 16
rect 5 3 9 6
rect 26 3 30 6
rect -2 2 34 3
rect 2 -2 14 2
rect 18 -2 34 2
rect -2 -3 34 -2
<< m1p >>
rect 2 43 6 47
rect 26 43 30 47
rect 10 33 14 37
rect 26 23 30 27
<< labels >>
rlabel metal1 4 0 4 0 4 gnd
rlabel metal1 4 100 4 100 4 vdd
rlabel metal1 4 45 4 45 4 A
rlabel metal1 12 35 12 35 4 B
rlabel metal1 28 45 28 45 4 Y
rlabel metal1 28 25 28 25 4 C
<< end >>
