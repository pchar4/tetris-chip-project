magic
tech scmos
timestamp 1711307567
<< metal1 >>
rect -10 2 10 3
rect 9 -2 10 2
rect -10 -3 10 -2
<< m2contact >>
rect -10 -2 9 2
<< metal2 >>
rect -10 2 10 3
rect 9 -2 10 2
rect -10 -3 10 -2
<< end >>
