/clear/apps/osu/soc-2.7/cadence/lib/ami05/lib/osu05_stdcells.lef