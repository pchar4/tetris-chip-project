// testbench just for the FSM

module fsm_tb();

reg in_clka, in_clkb, restart, touched, new_piece;
reg [3:0] which_row;
reg [1:0] state;

// creating an FSM


endmodule
