magic
tech scmos
timestamp 1712256841
<< nwell >>
rect -7 48 35 105
<< ntransistor >>
rect 7 6 9 16
rect 15 6 17 16
rect 23 6 25 26
<< ptransistor >>
rect 7 54 9 94
rect 12 54 14 94
rect 20 54 22 94
<< ndiffusion >>
rect 20 24 23 26
rect 18 22 23 24
rect 2 15 7 16
rect 6 6 7 15
rect 9 15 15 16
rect 9 6 10 15
rect 14 6 15 15
rect 17 8 18 16
rect 22 8 23 22
rect 17 6 23 8
rect 25 25 30 26
rect 25 6 26 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 54 7 93
rect 9 54 12 94
rect 14 93 20 94
rect 14 54 15 93
rect 19 54 20 93
rect 22 93 27 94
rect 22 54 23 93
<< ndcontact >>
rect 2 6 6 15
rect 10 6 14 15
rect 18 8 22 22
rect 26 6 30 25
<< pdcontact >>
rect 2 54 6 93
rect 15 54 19 93
rect 23 54 27 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 12 94 14 96
rect 20 94 22 96
rect 7 53 9 54
rect 6 51 9 53
rect 6 19 8 51
rect 12 41 14 54
rect 20 51 22 54
rect 20 49 25 51
rect 16 37 17 39
rect 6 17 9 19
rect 7 16 9 17
rect 15 16 17 37
rect 23 26 25 49
rect 7 4 9 6
rect 15 4 17 6
rect 23 4 25 6
<< polycontact >>
rect 2 19 6 23
rect 19 45 23 49
rect 12 37 16 41
<< metal1 >>
rect -2 102 34 103
rect 2 98 14 102
rect 18 98 34 102
rect -2 97 34 98
rect 2 93 6 94
rect 15 93 19 97
rect 23 93 27 94
rect 2 51 6 54
rect 2 49 22 51
rect 2 48 19 49
rect 27 47 30 57
rect 10 33 15 37
rect 20 30 23 45
rect 26 43 30 47
rect 11 27 23 30
rect 2 23 6 27
rect 11 16 14 27
rect 27 26 30 43
rect 26 25 30 26
rect 2 15 6 16
rect 10 15 14 16
rect 18 22 22 24
rect 2 3 6 6
rect 18 3 22 8
rect -2 2 34 3
rect 2 -2 14 2
rect 18 -2 34 2
rect -2 -3 34 -2
<< m1p >>
rect 26 43 30 47
rect 10 33 14 37
rect 2 23 6 27
<< labels >>
rlabel metal1 28 45 28 45 4 Y
rlabel metal1 12 35 12 35 4 B
rlabel metal1 4 100 4 100 4 vdd
rlabel metal1 4 0 4 0 4 gnd
rlabel metal1 4 25 4 25 4 A
<< end >>
