magic
tech scmos
timestamp 1712256841
<< m2contact >>
rect -2 -2 2 2
<< end >>
