magic
tech scmos
timestamp 1712020386
<< end >>
